CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 12 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
270 130 30 200 9
93 93 1333 746
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 Z:\home\matheussm\Documentos\UFCG\P1\IC\Circuit Maker\BOM.DAT
0 7
93 93 1333 746
143654930 0
0
6 Title:
5 Name:
0
0
0
7
13 Logic Switch~
5 423 315 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21088 0
2 5V
-6 -16 8 -8
1 C
-4 -16 3 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 424 278 0 1 11
0 5
0
0 0 21088 0
2 0V
-6 -16 8 -8
1 B
-2 -16 5 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 424 241 0 1 11
0 7
0
0 0 21088 0
2 0V
-6 -16 8 -8
1 A
-3 -17 4 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
14 Logic Display~
6 599 261 0 1 2
12 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
9 Inverter~
13 463 278 0 2 22
0 5 4
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
5394 0 0
0
0
9 Inverter~
13 466 239 0 2 22
0 7 6
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
7734 0 0
0
0
9 3-In AND~
219 545 277 0 4 22
0 6 4 3 2
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 AND
-16 -25 5 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 1 0
1 U
9914 0 0
0
0
6
4 1 2 0 0 8320 0 7 4 0 0 3
566 277
566 279
599 279
1 3 3 0 0 4224 0 1 7 0 0 5
435 315
505 315
505 296
521 296
521 286
2 2 4 0 0 8320 0 5 7 0 0 3
484 278
484 277
521 277
1 1 5 0 0 4224 0 2 5 0 0 2
436 278
448 278
2 1 6 0 0 8320 0 6 7 0 0 5
487 239
505 239
505 260
521 260
521 268
1 1 7 0 0 4224 0 3 6 0 0 3
436 241
451 241
451 239
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 39
433 170 602 214
437 172 598 204
39  QUEST�O 8(ITEM A)
SA�DA COM PORTA AND
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
