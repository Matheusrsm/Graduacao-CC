CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 10 9 100 9
0 66 640 394
7 5.000 V
7 5.000 V
3 GND
1.66667e+006 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 394
8912898 0
0
0
0
0
0
0
23
13 Logic Switch~
5 61 269 0 1 11
0 4
0
0 0 4448 0
2 5V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 60 220 0 1 11
0 5
0
0 0 4448 0
2 5V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 60 169 0 1 11
0 6
0
0 0 4448 0
2 5V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 59 120 0 1 11
0 7
0
0 0 4448 0
2 5V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
10 2-In NAND~
219 147 278 0 3 21
0 4 3 13
0
0 0 96 0
6 74LS00
-14 -24 28 -16
3 U1D
-4 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
5394 0 0
0
0
10 2-In NAND~
219 146 229 0 3 21
0 5 3 14
0
0 0 96 0
6 74LS00
-14 -24 28 -16
3 U1C
-4 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
7734 0 0
0
0
10 2-In NAND~
219 147 178 0 3 21
0 6 3 15
0
0 0 96 0
6 74LS00
-14 -24 28 -16
3 U1B
-4 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
9914 0 0
0
0
10 2-In NAND~
219 142 129 0 3 21
0 7 3 16
0
0 0 96 0
6 74LS00
-14 -24 28 -16
3 U1A
-4 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 2 0
1 U
3747 0 0
0
0
7 Ground~
168 74 86 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
11 Signal Gen~
195 35 50 0 24 64
0 3 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1232348160 0 1084227584
0 841731191 841731191 882970544 897988541
20
0 1e+006 0 5 0 1e-008 1e-008 3e-007 1e-006 0
0 0 0 0 0 0 0 0 0 0
0
0 0 320 0
4 0/5V
-14 -28 14 -20
2 V5
-7 -38 7 -30
0
0
42 %D %1 %2 DC 0 PULSE(0 5 0 10n 10n 300n 1u)
0
0
4 SIP3
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
2 +V
167 338 25 0 1 3
0 8
0
0 0 53600 0
4 +15V
9 -2 37 6
2 V6
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9325 0 0
0
0
7 Ground~
168 232 160 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
7 Ground~
168 300 210 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
7 Ground~
168 369 260 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
7 Ground~
168 438 307 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
12 NPN Trans:C~
219 227 129 0 3 7
0 12 16 2
12 NPN Trans:C~
0 0 320 0
3 NPN
17 -5 38 3
2 Q1
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
4718 0 0
0
0
12 NPN Trans:C~
219 295 178 0 3 7
0 11 15 2
12 NPN Trans:C~
0 0 320 0
3 NPN
17 -5 38 3
2 Q2
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
3874 0 0
0
0
12 NPN Trans:C~
219 364 229 0 3 7
0 10 14 2
12 NPN Trans:C~
0 0 320 0
3 NPN
17 -5 38 3
2 Q3
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
6671 0 0
0
0
12 NPN Trans:C~
219 433 278 0 3 7
0 9 13 2
12 NPN Trans:C~
0 0 320 0
3 NPN
17 -5 38 3
2 Q4
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
3789 0 0
0
0
9 Resistor~
219 232 68 0 4 5
0 12 8 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 300 69 0 4 5
0 11 8 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3750 0 0
0
0
9 Resistor~
219 369 69 0 4 5
0 10 8 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 438 70 0 4 5
0 9 8 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
538 0 0
0
0
25
2 0 3 0 0 4096 0 8 0 0 2 2
118 138
88 138
1 2 3 0 0 8320 0 10 5 0 0 4
66 45
88 45
88 287
123 287
2 1 2 0 0 8320 0 10 9 0 0 3
66 55
74 55
74 80
2 0 3 0 0 0 0 6 0 0 2 2
122 238
88 238
2 0 3 0 0 0 0 7 0 0 2 2
123 187
88 187
1 1 4 0 0 4224 0 1 5 0 0 2
73 269
123 269
1 1 5 0 0 4224 0 2 6 0 0 2
72 220
122 220
1 1 6 0 0 4224 0 3 7 0 0 2
72 169
123 169
1 1 7 0 0 4224 0 4 8 0 0 2
71 120
118 120
1 0 8 0 0 4096 0 11 0 0 13 2
338 34
338 43
2 0 8 0 0 12288 0 22 0 0 13 4
369 51
369 55
369 55
369 43
2 0 8 0 0 0 0 21 0 0 13 4
300 51
300 54
300 54
300 43
2 2 8 0 0 8320 0 20 23 0 0 4
232 50
232 43
438 43
438 52
3 1 2 0 0 0 0 19 15 0 0 2
438 296
438 301
3 1 2 0 0 0 0 18 14 0 0 2
369 247
369 254
3 1 2 0 0 0 0 17 13 0 0 2
300 196
300 204
3 1 2 0 0 0 0 16 12 0 0 2
232 147
232 154
1 1 9 0 0 4224 0 23 19 0 0 2
438 88
438 260
1 1 10 0 0 4224 0 22 18 0 0 2
369 87
369 211
1 1 11 0 0 4224 0 21 17 0 0 2
300 87
300 160
1 1 12 0 0 4224 0 20 16 0 0 2
232 86
232 111
3 2 13 0 0 4224 0 5 19 0 0 2
174 278
415 278
3 2 14 0 0 4224 0 6 18 0 0 2
173 229
346 229
3 2 15 0 0 4224 0 7 17 0 0 2
174 178
277 178
3 2 16 0 0 4224 0 8 16 0 0 2
169 129
209 129
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 3e-006 2.5e-008 2.5e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1172 8534080 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
4.49983e-315 0 5.36094e-315 0 4.49983e-315 4.49983e-315
1040 0
4 1e-006 10
1
98 138
0 3 0 0 1	0 1 0 0
13352 8550464 100 100 0 0
77 66 977 276
4 417 1020 764
977 66
77 66
977 67
977 276
0 0
4.80844e-315 0 5.27183e-315 1.58818e-314 4.80864e-315 4.80864e-315
16 0
4 1e-006 10
1
300 68
0 11 0 0 1	0 20 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
