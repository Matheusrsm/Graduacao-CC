CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 3
0 66 640 343
7 5.000 V
7 5.000 V
3 GND
0 343 640 452
16777218 0
0
1  
1  
1  
1  
1  
17
13 Logic Switch~
5 38 51 0 2 3
0 15 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 S1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 37 70 0 2 3
0 14 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 S2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 177 30 0 2 3
0 17 -99
0
0 0 20592 0
2 5V
-7 -16 7 -8
2 S3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 177 10 0 2 3
0 16 -99
0
0 0 20592 0
2 5V
-7 -16 7 -8
2 S4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 147 195 0 2 3
0 9 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 S5
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
12 Hex Display~
7 319 153 0 4 9
10 5 6 7 2
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -52 17 -44
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7734 0 0
0
0
12 Hex Display~
7 241 42 0 4 9
10 10 11 12 13
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -52 17 -44
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9914 0 0
0
0
14 Logic Display~
6 248 167 0 1 3
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
9 2-In AND~
219 214 219 0 3 21
0 9 8 3
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U2A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 3 0
1 U
3549 0 0
0
0
9 Inverter~
13 130 228 0 2 21
0 4 8
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 4 1 0
1 U
7931 0 0
0
0
5 SCOPE
12 446 141 0 3 3
0 7 -99 65
0
0 0 61680 0
2 A3
-7 -4 7 4
2 V1
-7 -14 7 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
5 SCOPE
12 409 141 0 3 3
0 6 -99 65
0
0 0 61680 0
2 A2
-7 -4 7 4
2 V2
-7 -14 7 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
5 SCOPE
12 372 141 0 3 3
0 5 -99 65
0
0 0 61680 0
2 A1
-7 -4 7 4
2 V3
-7 -14 7 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
7 Ground~
168 310 245 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
7 Pulser~
4 40 111 0 9 9
0 31 32 4 33 -99 0 5 5 4
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7668 0 0
0
0
7 74LS168
8 132 97 0 14 29
0 15 14 4 34 35 36 37 17 16
38 13 12 11 10
0
0 0 12528 0
8 74LS168A
-28 -60 28 -52
2 U3
-7 -70 7 -62
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 -33686019
65 0 0 512 1 1 0 0
1 U
4718 0 0
0
0
5 Macro
94 398 221 0 3 7
0 5 6 7
5 Macro
1 0 4240 0
0
0
0
0
0
0
0
0
7

0 0 0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3874 0 0
0
0
20
1 3 3 0 0 4224 0 8 9 0 0 3
248 185
248 219
235 219
1 0 4 0 0 8320 0 10 0 0 12 3
115 228
82 228
82 102
1 1 5 0 0 4096 0 17 6 0 0 3
366 212
328 212
328 177
2 2 6 0 0 4096 0 17 6 0 0 3
366 221
322 221
322 177
3 3 7 0 0 8320 0 17 6 0 0 4
430 221
430 236
316 236
316 177
1 0 7 0 0 0 0 11 0 0 5 3
446 153
446 236
430 236
1 0 6 0 0 8320 0 12 0 0 4 4
409 153
409 177
353 177
353 221
1 0 5 0 0 12416 0 13 0 0 3 4
372 153
372 169
345 169
345 212
4 1 2 0 0 4224 0 6 14 0 0 2
310 177
310 239
2 2 8 0 0 4224 0 10 9 0 0 2
151 228
190 228
1 1 9 0 0 12416 0 9 5 0 0 4
190 210
176 210
176 195
159 195
3 3 4 0 0 0 0 16 15 0 0 4
100 79
82 79
82 102
64 102
1 14 10 0 0 8320 0 7 16 0 0 3
250 66
250 133
164 133
2 13 11 0 0 8320 0 7 16 0 0 3
244 66
244 124
164 124
3 12 12 0 0 8320 0 7 16 0 0 3
238 66
238 115
164 115
4 11 13 0 0 8320 0 7 16 0 0 3
232 66
232 106
164 106
1 2 14 0 0 4224 0 2 16 0 0 2
49 70
94 70
1 1 15 0 0 4224 0 1 16 0 0 4
50 51
85 51
85 61
94 61
9 1 16 0 0 8320 0 16 4 0 0 4
164 70
200 70
200 10
189 10
1 8 17 0 0 8320 0 3 16 0 0 4
189 30
193 30
193 61
170 61
2
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 14
127 154 174 193
131 158 175 193
14 Toggle
Switch
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 25
256 78 327 119
260 82 328 117
25 Probe Wire 
To the Left
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 100 100 0 0
98 66 278 156
0 0 0 0
278 66
98 66
278 66
278 156
0 0
0.04 0 2 -0.4 0.04 2.4
0 0
0 2 5
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
0.005 0 0.8 -0.4 0.005 0.005
16 0
0 0.001 100
0
0 0 100 100 0 0
98 66 294 126
0 0 0 0
294 66
98 66
294 66
294 126
0 0
19108.5 10 56 60.2 19098.5 19098.5
12387 0
0 5000 10000
0
0 0 100 100 0 0
77 66 293 126
0 0 0 0
293 66
77 66
293 66
293 126
0 0
1e+006 1 -3.55271e-015 -3.55271e-015 999999 999999
4211 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
