CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 320 452
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 320 452
9961472 0
0
0
0
0
0
0
10
2 +V
167 204 167 0 1 64
0 4
0
0 0 54112 180
4 -15V
-13 11 15 19
3 VEE
-8 1 13 9
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
2 +V
167 204 92 0 1 64
0 5
0
0 0 54112 0
3 15V
-9 -16 12 -8
3 VCC
-8 -25 13 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
7 Ground~
168 131 206 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
11 Signal Gen~
195 38 124 0 24 64
0 8 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 1065353216 1148846080 -1082130432 1065353216
0 869711765 869711765 973279855 981668463
20
1 1000 -1 1 0 1e-007 1e-007 0.0005 0.001 0
0 0 0 0 0 0 0 0 0 0
0
0 0 576 0
5 -1/1V
-15 -48 20 -40
3 Vin
-11 -31 10 -23
0
0
52 %D %1 %2 DC 0 PULSE(-1 1 0 100n 100n 500u 1m) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
10 Polar Cap~
219 158 32 0 2 64
0 7 6
10 Polar Cap~
0 0 832 0
5 .02uf
-19 -18 16 -10
2 C2
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
10 Polar Cap~
219 155 119 0 2 64
0 7 3
10 Polar Cap~
0 0 832 0
5 .02uf
-19 -18 16 -10
2 C1
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
8 Op-Amp5~
219 204 125 0 5 64
0 2 3 5 4 6
8 Op-Amp5~
0 0 832 0
5 UA741
6 -16 41 -8
3 IC1
12 -27 33 -19
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 -33686019
88 0 0 256 1 1 0 0
1 U
9914 0 0
0
0
9 Resistor~
219 100 119 0 2 64
0 8 7
9 Resistor~
0 0 4960 0
5 39.8k
-17 -12 18 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 214 59 0 2 64
0 3 6
9 Resistor~
0 0 4960 0
4 159k
-14 -12 14 -4
2 RF
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 131 153 0 3 64
0 2 7 -1
9 Resistor~
0 0 4960 90
5 401.9
5 1 40 9
2 R2
17 -10 31 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
13
1 0 3 0 0 8320 0 9 0 0 2 3
196 59
177 59
177 119
2 2 3 0 0 0 0 6 7 0 0 2
161 119
186 119
4 1 4 0 0 4224 0 7 1 0 0 2
204 138
204 152
1 3 5 0 0 4224 0 2 7 0 0 2
204 101
204 112
5 2 6 0 0 8192 0 7 9 0 0 4
222 125
253 125
253 59
232 59
1 0 2 0 0 4096 0 3 0 0 11 2
131 200
131 185
1 0 2 0 0 0 0 10 0 0 11 2
131 171
131 185
2 0 6 0 0 4224 0 5 0 0 5 3
164 32
253 32
253 59
0 1 7 0 0 4224 0 0 5 10 0 3
131 119
131 32
147 32
2 0 7 0 0 0 0 10 0 0 13 2
131 135
131 119
2 1 2 0 0 12416 0 4 7 0 0 6
69 129
71 129
71 185
178 185
178 131
186 131
1 1 8 0 0 4224 0 8 4 0 0 2
82 119
69 119
1 2 7 0 0 0 0 6 8 0 0 2
144 119
118 119
0
0
25 0 0
0
0
0
0 0 0
0
0 0 0
100 0 1 2000
0 0.005 2.5e-005 2.5e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3704 8519744 100 100 0 0
77 66 287 126
320 66 640 259
287 66
77 66
287 66
287 126
0 0
0 0 0 0 0 0
16 0
4 0.001 10
2
76 119
0 8 0 0 1	0 12 0 0
253 105
0 6 0 0 2	0 5 0 0
2752 1472576 100 100 0 0
77 66 287 126
0 66 140 136
287 66
77 66
287 66
287 126
0 0
0 0 0 0 0 0
16 0
4 5e-006 10
1
204 107
0 5 0 0 1	0 4 0 0
2840 4356160 100 100 0 0
77 66 287 126
320 259 640 452
287 66
77 66
287 67
287 126
0 0
0 0 0 0 0 0
16 0
4 500 1000
1
253 112
0 6 0 0 2	0 5 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
