CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 640 452
7 5.000 V
7 5.000 V
3 GND
0 66 640 452
9437184 0
0
0
0
0
0
0
14
9 Inverter~
13 346 224 0 2 21
0 6 17
0
0 0 112 90
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 1 1 0
1 U
8953 0 0
0
0
13 Piezo Buzzer~
174 481 213 0 2 5
10 4 2
0
0 0 4208 0
4 .1uF
10 -16 38 -8
0
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
2 BZ
4441 0 0
0
0
14 Logic Display~
6 509 79 0 1 3
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
6 74LS74
17 403 208 0 12 25
0 35 36 17 16 37 38 39 40 4
41 42 43
0
0 0 12464 0
6 74LS74
-21 -60 21 -52
0
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 -33686019
65 0 0 512 1 1 0 0
1 U
6153 0 0
0
0
14 NO PushButton~
191 472 120 0 2 5
0 2 15
0
0 0 20592 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5394 0 0
0
0
14 NO PushButton~
191 375 120 0 2 5
0 2 16
0
0 0 20592 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7734 0 0
0
0
7 Window~
179 270 212 0 4 9
0 6 5 44 45
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 WND
9914 0 0
0
0
8 Hex Key~
166 227 40 0 11 11
0 7 8 9 10 0 0 0 0 0
0 48
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3747 0 0
0
0
8 Hex Key~
166 190 40 0 11 11
0 11 12 13 14 0 0 0 0 0
4 52
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3549 0 0
0
0
7 Ground~
168 519 276 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
7 Window~
179 146 217 0 4 9
0 6 5 46 47
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 WND
9325 0 0
0
0
7 Window~
179 37 218 0 4 9
0 6 5 48 49
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 WND
8903 0 0
0
0
5 Delay
94 280 101 0 11 23
0 14 13 12 11 10 9 8 7 5
15 16
5 Delay
1 0 4240 0
0
0
0
0
0
0
0
0
23

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
9 Resistor~
219 473 261 0 4 5
0 6 2 0 -1
9 Resistor~
0 0 4208 0
2 1k
-7 -12 7 -4
0
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3363 0 0
0
0
25
2 0 2 0 0 4096 0 2 0 0 7 2
512 213
519 213
9 1 4 0 0 8320 0 4 2 0 0 4
435 181
445 181
445 213
450 213
0 1 5 0 0 4096 0 0 3 21 0 3
326 152
509 152
509 97
1 1 6 0 0 12416 0 12 14 0 0 4
83 236
89 236
89 261
455 261
1 0 2 0 0 12288 0 6 0 0 7 4
392 128
413 128
413 144
519 144
2 0 2 0 0 0 0 14 0 0 7 2
491 261
519 261
1 1 2 0 0 8320 0 5 10 0 0 3
489 128
519 128
519 270
1 0 6 0 0 0 0 11 0 0 4 3
192 235
205 235
205 261
2 0 5 0 0 0 0 11 0 0 21 3
192 226
206 226
206 163
8 1 7 0 0 8320 0 13 8 0 0 3
248 137
236 137
236 64
2 7 8 0 0 4224 0 8 13 0 0 3
230 64
230 128
248 128
3 6 9 0 0 4224 0 8 13 0 0 3
224 64
224 119
248 119
5 4 10 0 0 8320 0 13 8 0 0 3
248 110
218 110
218 64
1 4 11 0 0 8320 0 9 13 0 0 3
199 64
199 101
248 101
2 3 12 0 0 8320 0 9 13 0 0 3
193 64
193 92
248 92
3 2 13 0 0 8320 0 9 13 0 0 3
187 64
187 83
248 83
1 4 14 0 0 4224 0 13 9 0 0 3
248 74
181 74
181 64
10 2 15 0 0 4224 0 13 5 0 0 4
318 137
429 137
429 128
455 128
4 0 16 0 0 8320 0 4 0 0 20 3
365 199
338 199
338 128
11 2 16 0 0 0 0 13 6 0 0 2
318 128
358 128
9 2 5 0 0 12416 0 13 12 0 0 6
312 83
326 83
326 163
89 163
89 227
83 227
2 3 17 0 0 4224 0 1 4 0 0 3
349 206
349 190
365 190
1 0 6 0 0 0 0 1 0 0 4 2
349 242
349 261
1 0 6 0 0 0 0 7 0 0 4 3
316 230
326 230
326 261
2 0 5 0 0 0 0 7 0 0 21 3
316 221
326 221
326 163
4
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 18
247 12 336 62
251 16 326 54
18 Exit Delay 
Time
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 13
440 57 507 107
444 61 497 99
13 Enable
Alarm
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 12
350 57 417 107
354 61 407 99
12 Reset
Alarm
-19 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 91
10 24 220 164
14 28 208 138
91 Normally-Open
Parallel Circuit
Burgler Alarm
With Latched Alarm 
Signal And Exit Delay
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 100 100 0 0
77 66 617 126
0 0 0 0
617 66
77 66
617 66
617 126
0 0
0.0005 0 1.2 -1.2 0.0005 0.0005
16 0
0 0.0001 10
0
0 0 100 100 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 -1.#IND -1.#IND 0 0
0 0
0 0.0002 10
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
