CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 80 9
0 66 640 343
7 5.000 V
7 5.000 V
3 GND
100000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 343
11010054 0
0
0
0
0
0
0
36
13 Logic Switch~
5 154 271 0 1 11
0 4
0
0 0 4448 0
2 0V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 156 298 0 1 11
0 5
0
0 0 4448 0
2 0V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
5 SAVE-
218 246 254 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 C
3 -26 10 -18
5 SAVE1
-11 -36 24 -28
0
0
11 *TRAN 0 5 0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 1 0 0 0
4 SAVE
3618 0 0
0
0
9 Inverter~
13 568 324 0 2 21
0 9 15
0
0 0 96 0
4 4069
-14 -19 14 -11
3 U4B
-11 -29 10 -21
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 2 4 0
1 U
6153 0 0
0
0
9 Inverter~
13 569 274 0 2 21
0 10 14
0
0 0 96 0
4 4069
-14 -19 14 -11
3 U4A
-11 -29 10 -21
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 1 4 0
1 U
5394 0 0
0
0
9 Inverter~
13 568 230 0 2 21
0 16 13
0
0 0 96 0
4 4069
-14 -19 14 -11
3 U1F
-11 -29 10 -21
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 6 1 0
1 U
7734 0 0
0
0
9 Inverter~
13 568 186 0 2 21
0 6 12
0
0 0 96 0
4 4069
-14 -19 14 -11
3 U1E
-11 -29 10 -21
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 5 1 0
1 U
9914 0 0
0
0
10 2-In NAND~
219 213 285 0 3 21
0 4 5 11
0
0 0 96 0
6 74LS00
-14 -24 28 -16
3 U6A
-4 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 6 0
1 U
3747 0 0
0
0
6 74112~
219 506 160 0 7 31
0 8 8 10 8 11 25 9
0
0 0 4192 0
7 74LS112
-3 -60 46 -52
3 U3A
11 -70 32 -62
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -33686019
65 0 0 512 2 1 3 0
1 U
3549 0 0
0
0
6 74112~
219 418 160 0 7 31
0 8 8 16 8 11 26 10
0
0 0 4192 0
7 74LS112
-3 -60 46 -52
3 U2A
11 -70 32 -62
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -33686019
65 0 0 512 2 1 2 0
1 U
7931 0 0
0
0
6 74112~
219 327 159 0 7 31
0 8 8 6 8 11 27 16
0
0 0 4192 0
7 74LS112
-3 -60 46 -52
3 U5B
11 -70 32 -62
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -33686019
65 0 0 512 2 2 5 0
1 U
9325 0 0
0
0
6 74112~
219 245 158 0 7 31
0 8 8 3 8 11 28 6
0
0 0 4192 0
7 74LS112
-3 -60 46 -52
3 U5A
11 -70 32 -62
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -33686019
65 0 0 512 2 1 5 0
1 U
8903 0 0
0
0
5 SAVE-
218 302 186 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
11 *TRAN 0 5 0
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
5 SAVE-
218 200 165 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
11 *TRAN 0 5 0
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
3363 0 0
0
0
2 +V
167 698 66 0 1 3
0 7
0
0 0 53600 0
4 +15V
-14 -22 14 -14
2 V3
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7668 0 0
0
0
7 Ground~
168 765 363 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4718 0 0
0
0
7 Ground~
168 721 308 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3874 0 0
0
0
7 Ground~
168 675 261 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
7 Ground~
168 619 215 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3789 0 0
0
0
2 +V
167 340 64 0 1 3
0 8
0
0 0 53600 0
3 +5V
-10 -15 11 -7
2 V4
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4871 0 0
0
0
12 NPN Trans:C~
219 614 186 0 3 7
0 20 12 2
12 NPN Trans:C~
0 0 320 0
3 NPN
17 -5 38 3
2 Q1
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
3750 0 0
0
0
12 NPN Trans:C~
219 670 230 0 3 7
0 19 13 2
12 NPN Trans:C~
0 0 320 0
3 NPN
17 -5 38 3
2 Q2
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
8778 0 0
0
0
12 NPN Trans:C~
219 716 274 0 3 7
0 18 14 2
12 NPN Trans:C~
0 0 320 0
3 NPN
17 -5 38 3
2 Q3
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
538 0 0
0
0
12 NPN Trans:C~
219 760 324 0 3 7
0 17 15 2
12 NPN Trans:C~
0 0 320 0
3 NPN
17 -5 38 3
2 Q4
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
6843 0 0
0
0
4 .IC~
207 24 169 0 1 3
0 23
0
0 0 53568 0
2 0V
-7 -15 7 -7
4 CMD1
-14 -25 14 -17
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
3 CMD
3136 0 0
0
0
2 +V
167 103 78 0 1 3
0 21
0
0 0 53600 0
3 +5V
-11 -22 10 -14
2 V5
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5950 0 0
0
0
10 555 Timer~
219 141 143 0 8 17
0 2 23 3 21 22 23 24 21
10 555 Timer~
0 0 6464 0
3 555
-10 -23 11 -15
2 U7
-7 -33 7 -25
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 -33686019
88 0 0 0 1 1 0 0
1 U
5670 0 0
0
0
10 Polar Cap~
219 52 218 0 2 5
0 23 2
10 Polar Cap~
0 0 832 26894
5 .01uF
-48 2 -13 10
2 C1
-33 -8 -19 0
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
6828 0 0
0
0
10 Polar Cap~
219 176 213 0 2 5
0 22 2
10 Polar Cap~
0 0 832 26894
5 .01uF
10 4 45 12
2 C2
21 -6 35 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
6735 0 0
0
0
7 Ground~
168 90 252 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8365 0 0
0
0
9 Resistor~
219 619 134 0 4 5
0 20 7 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 675 137 0 4 5
0 19 7 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
4551 0 0
0
0
9 Resistor~
219 721 137 0 4 5
0 18 7 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3635 0 0
0
0
9 Resistor~
219 765 140 0 4 5
0 17 7 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3973 0 0
0
0
9 Resistor~
219 51 173 0 2 5
0 23 24
9 Resistor~
0 0 4960 90
3 500
4 0 25 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3851 0 0
0
0
9 Resistor~
219 51 116 0 4 5
0 24 21 0 1
9 Resistor~
0 0 4960 90
3 100
7 0 28 8
2 R6
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
8383 0 0
0
0
55
0 1 2 0 0 4096 0 0 30 46 0 4
90 235
90 248
90 248
90 246
3 3 3 0 0 12416 0 27 12 0 0 6
109 152
98 152
98 179
200 179
200 131
215 131
1 1 4 0 0 4224 0 1 8 0 0 4
166 271
179 271
179 276
189 276
1 2 5 0 0 12416 0 2 8 0 0 4
168 298
178 298
178 294
189 294
3 0 6 0 0 4096 0 11 0 0 6 2
297 132
283 132
7 1 6 0 0 12416 0 12 7 0 0 4
269 122
283 122
283 186
553 186
1 0 7 0 0 4096 0 15 0 0 36 2
698 75
698 99
1 0 8 0 0 4096 0 11 0 0 21 2
327 96
327 84
7 1 9 0 0 8320 0 9 4 0 0 4
530 124
543 124
543 324
553 324
0 1 10 0 0 4224 0 0 5 22 0 3
455 133
455 274
554 274
1 0 8 0 0 8192 0 9 0 0 21 3
506 97
506 84
464 84
1 0 8 0 0 0 0 10 0 0 21 2
418 97
418 84
1 0 8 0 0 0 0 12 0 0 21 2
245 95
245 84
1 0 8 0 0 0 0 20 0 0 21 2
340 73
340 84
2 0 8 0 0 0 0 9 0 0 21 2
482 124
464 124
2 0 8 0 0 0 0 10 0 0 17 2
394 124
378 124
4 0 8 0 0 8192 0 10 0 0 21 3
394 142
378 142
378 84
2 0 8 0 0 0 0 11 0 0 19 2
303 123
293 123
4 0 8 0 0 0 0 11 0 0 21 3
303 141
293 141
293 84
2 0 8 0 0 0 0 12 0 0 21 2
221 122
210 122
4 4 8 0 0 12416 0 12 9 0 0 6
221 140
210 140
210 84
464 84
464 142
482 142
7 3 10 0 0 0 0 10 9 0 0 4
442 124
455 124
455 133
476 133
5 0 11 0 0 4096 0 10 0 0 43 2
418 172
418 206
5 0 11 0 0 4096 0 11 0 0 43 2
327 171
327 206
2 2 12 0 0 4224 0 21 7 0 0 2
596 186
589 186
2 2 13 0 0 4224 0 6 22 0 0 2
589 230
652 230
2 2 14 0 0 4224 0 23 5 0 0 2
698 274
590 274
2 2 15 0 0 4224 0 4 24 0 0 2
589 324
742 324
1 0 16 0 0 4224 0 6 0 0 41 3
553 230
368 230
368 133
3 1 2 0 0 4096 0 24 16 0 0 2
765 342
765 357
3 1 2 0 0 0 0 23 17 0 0 2
721 292
721 302
3 1 2 0 0 0 0 22 18 0 0 2
675 248
675 255
3 1 2 0 0 0 0 21 19 0 0 2
619 204
619 209
2 0 7 0 0 0 0 33 0 0 36 2
721 119
721 99
2 0 7 0 0 0 0 32 0 0 36 2
675 119
675 99
2 2 7 0 0 8320 0 31 34 0 0 4
619 116
619 99
765 99
765 122
1 1 17 0 0 4224 0 34 24 0 0 2
765 158
765 306
1 1 18 0 0 4224 0 33 23 0 0 2
721 155
721 256
1 1 19 0 0 4224 0 32 22 0 0 2
675 155
675 212
1 1 20 0 0 4224 0 31 21 0 0 2
619 152
619 168
7 3 16 0 0 0 0 11 10 0 0 4
351 123
368 123
368 133
388 133
5 0 11 0 0 4096 0 12 0 0 43 2
245 170
245 206
3 5 11 0 0 12416 0 8 9 0 0 5
240 285
245 285
245 206
506 206
506 172
8 1 21 0 0 8192 0 27 26 0 0 3
173 134
173 87
103 87
1 0 2 0 0 8192 0 27 0 0 46 3
109 134
76 134
76 235
2 2 2 0 0 8320 0 29 28 0 0 4
175 220
175 235
51 235
51 225
5 1 22 0 0 8320 0 27 29 0 0 3
173 161
175 161
175 203
1 0 23 0 0 8192 0 25 0 0 49 3
24 181
24 192
51 192
0 0 23 0 0 4096 0 0 0 52 55 2
51 192
91 192
2 1 21 0 0 0 0 36 26 0 0 3
51 98
51 87
103 87
7 0 24 0 0 12416 0 27 0 0 53 6
173 143
188 143
188 112
86 112
86 143
51 143
1 1 23 0 0 0 0 35 28 0 0 2
51 191
51 208
1 2 24 0 0 0 0 36 35 0 0 2
51 134
51 155
4 1 21 0 0 8320 0 27 26 0 0 3
109 161
103 161
103 87
2 6 23 0 0 12416 0 27 27 0 0 6
109 143
91 143
91 192
186 192
186 152
173 152
5
-20 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 40
171 22 660 57
175 26 655 53
40 Mixed-mode Binary Ripple Counter Circuit
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
519 303 543 327
523 307 539 323
2 Q3
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
519 251 544 275
523 255 539 271
2 Q2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
519 208 543 232
523 212 539 228
2 Q1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
519 164 544 188
523 168 539 184
2 Q0
33 .OPTIONS ITL4=100.0 TRTOL=3.000

16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-005 5e-008 5e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2492 8526400 100 100 0 0
98 66 608 126
0 259 640 452
608 66
98 66
608 66
608 126
0 0
0 0 0 0 0 0
12409 0
4 1e-005 10
1
619 161
0 20 0 0 1	0 40 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
