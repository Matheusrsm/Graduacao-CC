CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
430 40 30 200 9
63 134 1370 772
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
54 C:\Users\H�rcules\Desktop\Circuito Maker\CM60S\BOM.DAT
0 7
63 134 1370 772
143655186 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 528 167 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-10 15 4 23
1 A
-5 -23 2 -15
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 537 301 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-5 18 9 26
1 B
-2 -30 5 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
14 Logic Display~
6 859 275 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 857 157 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
9 Inverter~
13 587 302 0 2 22
0 2 7
0
0 0 96 0
6 74LS04
-21 -19 21 -11
2 A1
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 3 0
1 U
5394 0 0
0
0
9 Inverter~
13 587 166 0 2 22
0 3 6
0
0 0 96 0
6 74LS04
-21 -19 21 -11
2 A2
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 3 0
1 U
7734 0 0
0
0
10 2-In NAND~
219 731 293 0 3 22
0 5 7 4
0
0 0 96 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
9914 0 0
0
0
10 2-In NAND~
219 730 175 0 3 22
0 6 4 5
0
0 0 96 0
4 7400
-7 -24 21 -16
2 A3
0 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 -1766218101
65 0 0 0 4 1 2 0
1 U
3747 0 0
0
0
8
1 1 2 0 0 8320 0 2 5 0 0 3
549 301
549 302
572 302
1 1 3 0 0 8320 0 1 6 0 0 3
540 167
540 166
572 166
1 0 4 0 0 4096 0 3 0 0 8 2
859 293
815 293
1 0 5 0 0 8192 0 4 0 0 7 3
857 175
857 177
816 177
2 1 6 0 0 8320 0 6 8 0 0 2
608 166
706 166
2 2 7 0 0 4224 0 5 7 0 0 2
608 302
707 302
3 1 5 0 0 16528 0 8 7 0 0 7
757 175
757 177
816 177
816 226
702 226
702 284
707 284
3 2 4 0 0 12416 0 7 8 0 0 6
758 293
815 293
815 244
694 244
694 184
706 184
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-006 1e-007 1e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
