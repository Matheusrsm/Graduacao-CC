CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
10 10 5 50 9
0 66 640 343
7 5.000 V
7 5.000 V
3 GND
62500 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 343 640 452
161480706 0
0
0
0
0
0
0
26
9 Data Seq~
170 364 228 0 17 21
0 19 20 21 22 23 24 25 5 26
27 51 1 80 1 1 0 81
0
0 0 20576 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -54 10 -46
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
0
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
8953 0 0
0
0
AAAAAAAAAAAAABABABABABAAAAAAAAAAABABABABABAAAAAAAAAAABABABABABAAAAAAAAAAABABABAB
ABAAAAAAAAAAABABABABABAAAAAAAAAAABABABABABAAAAAAAAAAABABABABABAAAAAAAAAAABABABAB
AB
6 Input~
177 632 94 0 17 17
0 3 0 0 0 0 0 0 0 0
83 105 103 49 32 32 32 32
0
0 0 53344 0
0
2 T1
-7 -26 7 -18
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4441 0 0
0
0
7 Output~
178 158 24 0 17 17
0 3 0 0 0 0 0 0 0 0
83 105 103 49 32 32 32 32
0
0 0 53344 0
0
2 T2
-13 -26 1 -18
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3618 0 0
0
0
7 Output~
178 158 45 0 17 17
0 4 0 0 0 0 0 0 0 0
83 105 103 50 32 32 32 32
0
0 0 53344 0
0
2 T3
-13 -26 1 -18
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6153 0 0
0
0
6 Input~
177 291 24 0 17 17
0 3 0 0 0 0 0 0 0 0
83 105 103 49 32 32 32 32
0
0 0 53344 0
0
2 T4
-7 -26 7 -18
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5394 0 0
0
0
6 Input~
177 633 151 0 17 17
0 4 0 0 0 0 0 0 0 0
83 105 103 50 32 32 32 32
0
0 0 53344 0
0
2 T5
-7 -26 7 -18
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7734 0 0
0
0
6 Input~
177 291 45 0 17 17
0 4 0 0 0 0 0 0 0 0
83 105 103 50 32 32 32 32
0
0 0 53344 0
0
2 T6
-7 -26 7 -18
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9914 0 0
0
0
9 Inverter~
13 508 84 0 2 21
0 4 3
0
0 0 96 0
4 4069
-14 -19 14 -11
3 U1A
-11 -29 10 -21
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 1 7 0
1 U
3747 0 0
0
0
12 Quad D Flop~
47 404 133 0 9 19
0 3 11 10 28 4 7 8 29 5
0
0 0 4192 0
4 QDFF
-14 -44 14 -36
2 U5
-7 -54 7 -46
0
15 DVCC=16;DGND=8;
81 %D [%16bi %8bi %1i %2i %3i %4i %9i][%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 -33686019
65 0 0 512 1 1 0 0
1 U
3549 0 0
0
0
9 Inverter~
13 508 147 0 2 21
0 8 9
0
0 0 96 0
4 4069
-14 -19 14 -11
3 U1B
-11 -29 10 -21
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 2 7 0
1 U
7931 0 0
0
0
9 Inverter~
13 508 115 0 2 21
0 7 12
0
0 0 96 0
4 4069
-14 -19 14 -11
3 U1C
-11 -29 10 -21
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 3 7 0
1 U
9325 0 0
0
0
8 2-In OR~
219 324 179 0 3 21
0 14 13 10
0
0 0 96 0
6 74LS32
-21 -24 21 -16
3 U4C
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 3 10 0
1 U
8903 0 0
0
0
8 2-In OR~
219 246 170 0 3 21
0 17 16 14
0
0 0 96 0
6 74LS32
-21 -24 21 -16
3 U4B
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 2 10 0
1 U
3834 0 0
0
0
8 2-In OR~
219 245 115 0 3 21
0 6 18 11
0
0 0 96 0
6 74LS32
-21 -24 21 -16
3 U4A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 10 0
1 U
3363 0 0
0
0
9 2-In AND~
219 252 246 0 3 21
0 15 12 13
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U3B
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 2 9 0
1 U
7668 0 0
0
0
9 2-In AND~
219 124 237 0 3 21
0 3 8 15
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U3A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 9 0
1 U
4718 0 0
0
0
9 2-In AND~
219 124 199 0 3 21
0 7 4 16
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2D
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 4 8 0
1 U
3874 0 0
0
0
9 2-In AND~
219 124 161 0 3 21
0 7 9 17
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2C
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 3 8 0
1 U
6671 0 0
0
0
9 2-In AND~
219 124 124 0 3 21
0 4 8 18
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2B
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 2 8 0
1 U
3789 0 0
0
0
9 2-In AND~
219 124 87 0 3 21
0 3 9 6
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 8 0
1 U
4871 0 0
0
0
5 SCOPE
12 297 333 0 3 3
0 4 0 49
0
0 0 61664 0
3 TP3
-11 -4 10 4
3 TP1
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3750 0 0
0
0
5 SCOPE
12 262 333 0 3 3
0 7 0 50
0
0 0 61664 0
3 TP2
-11 -4 10 4
3 TP2
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8778 0 0
0
0
5 SCOPE
12 226 333 0 3 3
0 8 0 51
0
0 0 61664 0
3 TP1
-11 -4 10 4
3 TP3
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
538 0 0
0
0
7 Ground~
168 169 409 0 3 3
0 2 0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6843 0 0
0
0
12 Hex Display~
7 178 340 0 9 19
10 4 7 8 2 0 2 2 2 2
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -52 17 -44
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3136 0 0
0
0
8 Speaker~
175 694 124 0 2 5
10 3 4
0
0 0 4192 0
1 8
-3 -22 4 -14
5 SPKR1
-17 -32 18 -24
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
3 SPK
5950 0 0
0
0
36
9 8 5 0 0 4224 0 9 1 0 0 3
404 169
404 264
396 264
1 1 3 0 0 4096 0 2 26 0 0 3
666 94
686 94
686 108
2 1 4 0 0 8192 0 26 6 0 0 3
686 140
686 151
667 151
2 1 3 0 0 12416 0 8 5 0 0 4
529 84
546 84
546 24
325 24
3 1 6 0 0 12416 0 20 14 0 0 4
145 87
185 87
185 106
232 106
1 0 4 0 0 4096 0 7 0 0 29 3
325 45
443 45
443 84
1 1 3 0 0 0 0 3 16 0 0 4
118 24
17 24
17 228
100 228
1 0 4 0 0 0 0 21 0 0 15 3
297 345
297 397
187 397
1 0 7 0 0 8192 0 22 0 0 18 3
262 345
262 386
181 386
1 0 8 0 0 8192 0 23 0 0 19 3
226 345
226 377
174 377
4 1 2 0 0 4224 0 25 24 0 0 2
169 364
169 403
2 0 9 0 0 4096 0 18 0 0 25 2
100 170
42 170
2 0 4 0 0 0 0 17 0 0 15 2
100 208
29 208
1 0 4 0 0 0 0 19 0 0 15 2
100 115
29 115
1 1 4 0 0 12416 0 25 4 0 0 5
187 364
187 397
29 397
29 45
118 45
0 0 7 0 0 8320 0 0 0 22 18 3
474 115
474 307
77 307
1 0 7 0 0 0 0 17 0 0 18 2
100 190
77 190
1 2 7 0 0 0 0 18 25 0 0 5
100 152
77 152
77 386
181 386
181 364
0 3 8 0 0 4096 0 0 25 28 0 4
102 297
102 377
175 377
175 364
3 3 10 0 0 8320 0 12 9 0 0 4
357 179
368 179
368 127
380 127
3 2 11 0 0 4224 0 14 9 0 0 2
278 115
380 115
1 6 7 0 0 0 0 11 9 0 0 2
493 115
428 115
2 0 8 0 0 0 0 16 0 0 28 2
100 246
66 246
2 2 12 0 0 12416 0 11 15 0 0 6
529 115
545 115
545 275
215 275
215 255
228 255
2 2 9 0 0 12416 0 10 20 0 0 6
529 147
535 147
535 287
42 287
42 96
100 96
0 1 8 0 0 0 0 0 10 28 0 2
440 147
493 147
1 0 3 0 0 0 0 9 0 0 4 3
380 103
369 103
369 24
2 7 8 0 0 12416 0 19 9 0 0 6
100 133
66 133
66 297
440 297
440 127
428 127
5 1 4 0 0 0 0 9 8 0 0 4
428 103
443 103
443 84
493 84
1 0 3 0 0 0 0 20 0 0 7 2
100 78
17 78
3 2 13 0 0 8320 0 15 12 0 0 4
273 246
294 246
294 188
311 188
3 1 14 0 0 4224 0 13 12 0 0 2
279 170
311 170
3 1 15 0 0 4224 0 16 15 0 0 2
145 237
228 237
2 3 16 0 0 4224 0 13 17 0 0 4
233 179
182 179
182 199
145 199
3 1 17 0 0 4224 0 18 13 0 0 2
145 161
233 161
3 2 18 0 0 4224 0 19 14 0 0 2
145 124
232 124
1
-17 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 70
329 337 636 385
333 341 640 389
70 This is a simple state machine with 
state sequence 0,3,4,5,2,7,6,1.
21 .OPTIONS METHOD=GEAR

2065 0 1
0
0
3 Vin
-0.1 0.1 0.005
3 Vee
-15 0 1
100 0 1 1e+006
0 8e-005 3.2e-007 3.2e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1248 1210432 100 100 0 0
0 0 0 0
0 66 140 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
4 1 2
0
1268 8525888 100 100 0 0
77 66 617 126
0 259 640 452
437 66
77 66
617 66
617 126
0 0
0 0 0 0 0 0
1024 0
2 2e-005 5
3
226 367
0 9 0 21 1	0 10 0 0
262 372
0 8 0 0 1	0 9 0 0
297 375
0 5 0 -17 1	0 8 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
