CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 300 100 9
0 66 640 452
7 5.000 V
7 5.000 V
3 GND
10000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 452
9961490 0
0
0
0
0
0
0
19
4 .IC~
207 282 73 0 1 64
0 3
0
0 0 53568 0
2 5V
-7 -15 7 -7
4 CMD1
-14 -25 14 -17
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
3 CMD
8953 0 0
0
0
4 .IC~
207 44 71 0 1 64
0 4
0
0 0 53568 0
2 0V
-7 -15 7 -7
4 CMD2
-14 -25 14 -17
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
3 CMD
4441 0 0
0
0
5 SAVE-
218 244 130 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 D
3 -26 10 -18
0
0
0
12 *TRAN 748m 8
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SAVE-
218 136 143 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 C
3 -26 10 -18
0
0
0
16 *TRAN -5.63 1.49
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
5 SAVE-
218 170 144 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
15 *TRAN -5.75 1.5
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SAVE-
218 78 118 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
12 *TRAN 748m 8
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
7 Ground~
168 243 230 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
7 Ground~
168 77 231 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
2 +V
167 162 29 0 1 64
0 5
0
0 0 53600 0
3 +8V
-10 -16 11 -8
2 V1
-7 -26 7 -18
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3549 0 0
0
0
12 NPN Trans:C~
219 238 157 0 3 64
0 3 7 8
12 NPN Trans:C~
0 0 320 0
6 2N3904
20 -4 62 4
2 Q1
34 -14 48 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 0 0 0
1 Q
7931 0 0
0
0
12 NPN Trans:C~
219 86 157 0 3 64
0 4 6 9
12 NPN Trans:C~
0 0 320 512
6 2N3904
-70 -5 -28 3
2 Q2
-56 -15 -42 -7
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 0 0 0
1 Q
9325 0 0
0
0
10 Capacitor~
219 106 124 0 2 64
0 4 7
10 Capacitor~
0 0 320 0
5 618pF
-12 -20 23 -12
2 C1
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
8903 0 0
0
0
10 Capacitor~
219 217 124 0 2 64
0 6 3
10 Capacitor~
0 0 320 0
6 1.55nF
-22 -19 20 -11
2 C2
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3834 0 0
0
0
6 Diode~
219 77 201 0 2 64
0 9 2
6 Diode~
0 0 320 26894
5 1N914
13 -2 48 6
2 D1
23 -12 37 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
3363 0 0
0
0
6 Diode~
219 243 198 0 2 64
0 8 2
6 Diode~
0 0 320 26894
5 1N914
14 -2 49 6
2 D2
24 -12 38 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
7668 0 0
0
0
9 Resistor~
219 77 85 0 4 64
0 4 5 0 1
9 Resistor~
0 0 352 90
2 1k
7 -2 21 6
2 R1
7 -12 21 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 135 86 0 4 64
0 7 5 0 1
9 Resistor~
0 0 352 90
3 47k
6 -5 27 3
2 R2
9 -15 23 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 243 88 0 4 64
0 3 5 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R3
8 -15 22 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 189 85 0 4 64
0 6 5 0 1
9 Resistor~
0 0 352 90
3 47k
7 -2 28 6
2 R4
10 -12 24 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
18
1 0 3 0 0 8320 0 1 0 0 13 3
282 85
282 107
243 107
1 0 4 0 0 8192 0 2 0 0 18 3
44 83
44 109
77 109
1 0 5 0 0 4096 0 9 0 0 6 2
162 38
162 54
2 0 5 0 0 0 0 19 0 0 6 2
189 67
189 54
2 0 5 0 0 0 0 17 0 0 6 2
135 68
135 54
2 2 5 0 0 8320 0 16 18 0 0 4
77 67
77 54
243 54
243 70
2 0 3 0 0 0 0 13 0 0 13 2
226 124
243 124
1 0 6 0 0 4096 0 13 0 0 11 2
208 124
189 124
2 0 7 0 0 4096 0 12 0 0 12 2
115 124
135 124
1 0 4 0 0 0 0 12 0 0 18 2
97 124
77 124
1 2 6 0 0 16512 0 19 11 0 0 5
189 103
189 144
163 144
163 157
100 157
1 2 7 0 0 8320 0 17 10 0 0 5
135 104
135 151
189 151
189 157
220 157
1 1 3 0 0 0 0 18 10 0 0 2
243 106
243 139
2 1 2 0 0 4224 0 15 7 0 0 2
243 208
243 224
3 1 8 0 0 4224 0 10 15 0 0 2
243 175
243 188
2 1 2 0 0 0 0 14 8 0 0 2
77 211
77 225
3 1 9 0 0 4224 0 11 14 0 0 2
77 175
77 191
1 1 4 0 0 4224 0 16 11 0 0 2
77 103
77 139
2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 418
321 42 585 366
325 46 581 302
418 The initial condition (.IC) 
devices are placed in this 
circuit to give the SPICE 
simulator a starting point for 
the outputs.  This allows the 
simulation to begin more 
quickly.  Since the circuit is 
not exactly symetrical (the 
capacitors are not the same), 
SPICE could begin the 
oscillation, but it would take 
a few moments to get it 
started.

Remove the .IC devices and try 
it!
-16 0 0 0 700 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 42
321 0 551 53
325 4 545 42
42 Collector Coupled 
Astable Multivibrator
0
16 0 1
0
0
0
0 0 0
0
0 0 0
200 0 1 1e+006
0 0.0005 1e-006 1e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
