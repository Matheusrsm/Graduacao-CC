CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 12 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
60 30 30 200 9
34 91 1332 708
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
53 C:\Users\Josefa Ramos\Documents\Circuit Maker\BOM.DAT
0 7
34 91 1332 708
143654930 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 178 221 0 1 11
0 3
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 S
-3 -18 4 -10
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 179 184 0 1 11
0 4
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 V
-2 -18 5 -10
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 180 150 0 1 11
0 5
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 D
-3 -17 4 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
14 Logic Display~
6 580 185 0 1 2
12 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
8 3-In OR~
219 517 203 0 4 22
0 8 7 6 2
0
0 0 624 0
4 4075
-14 -24 14 -16
2 OR
0 -25 14 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 2 0
1 U
5394 0 0
0
0
9 2-In AND~
219 368 267 0 3 22
0 4 3 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7734 0 0
0
0
9 2-In AND~
219 369 203 0 3 22
0 5 3 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9914 0 0
0
0
9 2-In AND~
219 369 138 0 3 22
0 5 4 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3747 0 0
0
0
10
4 1 2 0 0 4224 0 5 4 0 0 2
550 203
580 203
0 2 3 0 0 8320 0 0 6 4 0 3
212 221
212 276
344 276
0 1 4 0 0 8320 0 0 6 6 0 3
228 184
228 258
344 258
1 2 3 0 0 0 0 1 7 0 0 4
190 221
289 221
289 212
345 212
0 1 5 0 0 8320 0 0 7 7 0 3
211 150
211 194
345 194
1 2 4 0 0 0 0 2 8 0 0 4
191 184
253 184
253 147
345 147
1 1 5 0 0 0 0 3 8 0 0 4
192 150
244 150
244 129
345 129
3 3 6 0 0 12416 0 6 5 0 0 4
389 267
444 267
444 212
504 212
3 2 7 0 0 4224 0 7 5 0 0 2
390 203
505 203
3 1 8 0 0 12416 0 8 5 0 0 4
390 138
444 138
444 194
504 194
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 53
244 65 476 109
249 69 473 101
53 ITEM A - DIRETORIA DA ESCOLA
     SA�DA COM PORTA OR
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
