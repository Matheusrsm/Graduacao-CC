CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 800 319
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 800 319
10027026 1
0
6 Title:
5 Name:
0
0
0
10
2 +V
167 211 43 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
7 Ground~
168 119 147 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
5 SAVE-
218 330 123 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 G
3 -26 10 -18
0
0
0
30 *Combine
*TRAN 0.000 42.00 36
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3618 0 0
0
0
5 SAVE-
218 316 112 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 F
3 -26 10 -18
0
0
0
30 *Combine
*TRAN 0.000 42.00 30
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
6153 0 0
0
0
5 SAVE-
218 309 103 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 E
3 -26 10 -18
0
0
0
30 *Combine
*TRAN 0.000 42.00 24
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
5394 0 0
0
0
5 SAVE-
218 292 96 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 D
3 -26 10 -18
0
0
0
30 *Combine
*TRAN 0.000 42.00 18
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
7734 0 0
0
0
5 SAVE-
218 175 145 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
29 *Combine
*TRAN 0.000 42.00 6
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
9914 0 0
0
0
11 Signal Gen~
195 74 73 0 24 64
0 4 2 1 86 9 10 0 0 0
0 0 0 0 0 0 0 1145065161 0 1076090634
0 983730047 897988541 897988541 984245443
20
0 769.231 0 2.56 0 0.00124 1e-006 1e-006 0.0013 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 0/2.56V
-25 -30 24 -22
2 V4
-7 -40 7 -32
0
0
46 %D %1 %2 DC 0 PULSE(0 2.56 0 1.24m 1u 1u 1.3m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
2 +V
167 163 41 0 1 3
0 5
0
0 0 54128 0
5 2.56V
-17 -12 18 -4
2 V2
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3549 0 0
0
0
4 ADC8
219 253 86 0 14 29
0 4 5 2 10 3 10 9 8 7
6 11 12 13 14
4 ADC8
0 0 13040 0
4 ADC8
-14 -56 14 -48
2 U1
-7 -66 7 -58
0
15 DVCC=16;DGND=8;
98 %D [%16bi %8bi %1i %2i %3i %4i %5i]
+ [%16bo %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 -33686019
65 0 0 512 1 1 0 0
1 U
7931 0 0
0
0
10
1 5 3 0 0 4224 0 1 10 0 0 3
211 52
211 122
220 122
1 1 4 0 0 4224 0 8 10 0 0 2
105 68
220 68
3 0 2 0 0 4224 0 10 0 0 4 2
220 95
119 95
2 1 2 0 0 128 0 8 2 0 0 3
105 78
119 78
119 141
1 2 5 0 0 8320 0 9 10 0 0 3
163 50
163 86
220 86
10 0 6 0 0 4224 0 10 0 0 0 2
286 95
357 95
9 0 7 0 0 4224 0 10 0 0 0 2
286 104
357 104
8 0 8 0 0 4224 0 10 0 0 0 2
286 113
356 113
0 7 9 0 0 4224 0 0 10 0 0 2
361 122
286 122
6 4 10 0 0 12416 0 10 10 0 0 6
286 131
324 131
324 145
163 145
163 113
220 113
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-005 5e-007 5e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1724 8550464 100 100 0 0
77 66 767 186
0 319 800 572
113 66
96 66
767 126
767 126
0 0
3.13043e-006 1.65217e-006 0 0 5e-005 5e-005
13425 0
2 1e-005 5
5
309 122
0 9 0 37 1	0 9 0 0
312 113
0 8 0 15 1	0 8 0 0
313 104
0 7 0 -8 1	0 7 0 0
313 95
0 6 0 -32 1	0 6 0 0
186 145
0 10 0 -59 3	0 10 0 0
3420 8550464 100 100 0 0
77 66 977 246
0 403 1024 740
131 66
77 66
977 140
977 156
0 0
0.0002 0 0 0 0.0002 0.0002
13425 0
2 5e-005 10
8
199 103
0 12 0 -72 1	0 11 0 0
203 94
0 13 0 -50 1	0 11 0 0
203 85
0 14 0 -29 1	0 11 0 0
206 76
0 15 0 -10 1	0 11 0 0
325 85
0 11 0 16 1	0 11 0 0
330 94
0 10 0 35 1	0 11 0 0
334 112
0 9 0 55 1	0 11 0 0
339 121
0 8 0 71 1	0 11 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
