CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 800 319
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 800 319
10027026 1
0
6 Title:
5 Name:
0
0
0
18
5 SAVE-
218 317 121 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 G
3 -26 10 -18
5 SAVE1
-11 -36 24 -28
0
0
30 *Combine
*TRAN 0.000 42.00 36
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
8953 0 0
0
0
5 SAVE-
218 316 112 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 F
3 -26 10 -18
5 SAVE2
-11 -36 24 -28
0
0
30 *Combine
*TRAN 0.000 42.00 30
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
4441 0 0
0
0
5 SAVE-
218 316 94 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 E
3 -26 10 -18
5 SAVE3
-11 -36 24 -28
0
0
30 *Combine
*TRAN 0.000 42.00 24
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3618 0 0
0
0
5 SAVE-
218 315 85 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 D
3 -26 10 -18
5 SAVE4
-11 -36 24 -28
0
0
30 *Combine
*TRAN 0.000 42.00 18
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
6153 0 0
0
0
5 SAVE-
218 219 148 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 C
3 -26 10 -18
5 SAVE5
-11 -36 24 -28
0
0
30 *Combine
*TRAN 0.000 42.00 12
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
5394 0 0
0
0
5 SAVE-
218 223 122 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
5 SAVE6
-11 -36 24 -28
0
0
29 *Combine
*TRAN 0.000 42.00 6
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
7734 0 0
0
0
5 SAVE-
218 315 139 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
5 SAVE7
-11 -36 24 -28
0
0
29 *Combine
*TRAN 0.000 42.00 0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
9914 0 0
0
0
2 +V
167 162 55 0 1 3
0 3
0
0 0 54128 0
3 -12
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
11 Signal Gen~
195 392 164 0 24 64
0 6 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1232348160 0 1084227584
0 814313567 814313567 889599933 897988541
20
0 1e+006 0 5 0 1e-009 1e-009 5e-007 1e-006 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 512
4 0/5V
-9 -30 19 -22
2 V2
-2 -40 12 -32
0
0
40 %D %1 %2 DC 0 PULSE(0 5 0 1n 1n 500n 1u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3549 0 0
0
0
7 Ground~
168 117 199 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
7 Ground~
168 451 197 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
11 Signal Gen~
195 488 135 0 24 64
0 8 2 1 86 9 10 0 0 0
0 0 0 0 0 0 0 1120021696 0 1076090634
0 1009239468 897988541 897988541 1009303893
20
0 97.0874 0 2.56 0 0.01024 1e-006 1e-006 0.0103 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 512
7 0/2.56V
-20 -30 29 -22
2 V3
-2 -40 12 -32
0
0
48 %D %1 %2 DC 0 PULSE(0 2.56 0 10.24m 1u 1u 10.3m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
11 Signal Gen~
195 71 126 0 24 64
0 5 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1187205120 0 1084227584
897988541 814313567 814313567 906377149 942130604
20
0 25000 0 5 1e-006 1e-009 1e-009 2e-006 4e-005 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/5V
-14 -30 14 -22
2 V4
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 PULSE(0 5 1u 1n 1n 2u 40u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3834 0 0
0
0
7 Ground~
168 226 198 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
2 +V
167 394 51 0 1 3
0 9
0
0 0 54128 0
5 2.56V
-18 -22 17 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7668 0 0
0
0
7 Ground~
168 333 197 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4718 0 0
0
0
2 +V
167 216 54 0 1 3
0 4
0
0 0 54128 0
1 5
-4 -22 3 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3874 0 0
0
0
7 ADC0800
219 274 103 0 18 37
0 17 16 15 14 2 5 4 3 7
4 6 8 10 11 9 12 13 2
8 ADC0800~
0 0 4976 0
7 ADC0800
-25 -56 24 -48
2 U1
-7 -66 7 -58
0
0
68 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %10 %11 %12 %13 %14 %15 %16 %17 %18 %S
0
0
5 DIP18
37

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 1
2 3 4 5 6 7 8 9 10 11
12 13 14 15 16 17 18 -1610612644
88 0 0 0 1 1 0 0
1 U
6671 0 0
0
0
21
1 8 3 0 0 8320 0 8 18 0 0 3
162 64
162 139
241 139
7 0 4 0 0 4096 0 18 0 0 5 2
241 130
216 130
2 0 2 0 0 4096 0 9 0 0 4 2
367 169
333 169
18 1 2 0 0 8320 0 18 16 0 0 3
307 76
333 76
333 191
1 10 4 0 0 4224 0 17 18 0 0 5
216 63
216 163
312 163
312 148
307 148
6 1 5 0 0 4224 0 18 13 0 0 2
241 121
102 121
1 11 6 0 0 12416 0 9 18 0 0 4
367 159
355 159
355 139
307 139
9 0 7 0 0 4224 0 18 0 0 0 2
241 148
183 148
12 1 8 0 0 4224 0 18 12 0 0 2
307 130
463 130
2 1 2 0 0 0 0 13 10 0 0 3
102 131
117 131
117 193
2 1 2 0 0 0 0 12 11 0 0 3
463 140
451 140
451 191
5 1 2 0 0 0 0 18 14 0 0 3
241 112
226 112
226 192
15 1 9 0 0 4224 0 18 15 0 0 3
307 103
394 103
394 60
13 0 10 0 0 4224 0 18 0 0 0 2
307 121
368 121
14 0 11 0 0 4224 0 18 0 0 0 2
307 112
367 112
16 0 12 0 0 4224 0 18 0 0 0 2
307 94
376 94
17 0 13 0 0 4224 0 18 0 0 0 2
307 85
374 85
4 0 14 0 0 4224 0 18 0 0 0 2
241 103
183 103
3 0 15 0 0 4224 0 18 0 0 0 2
241 94
184 94
2 0 16 0 0 4224 0 18 0 0 0 2
241 85
181 85
1 0 17 0 0 4224 0 18 0 0 0 2
241 76
181 76
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.0005 5e-007 5e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2032 8550464 100 100 0 0
77 66 767 186
0 319 800 572
163 66
77 66
767 142
767 126
0 0
2.24348e-005 0 -8 0 0.000193001 0.000193001
13425 0
2 3e-005 10
7
317 139
0 6 0 -59 3	0 7 0 0
132 121
0 5 0 -44 1	0 6 0 0
197 148
0 7 0 -27 1	0 8 0 0
313 121
0 10 0 -11 1	0 14 0 0
313 112
0 11 0 8 1	0 15 0 0
314 94
0 12 0 25 1	0 16 0 0
314 85
0 13 0 43 1	0 17 0 0
3420 8550464 100 100 0 0
77 66 977 246
0 403 1024 740
131 66
77 66
977 140
977 156
0 0
4.75121e-315 0 0 0 4.75121e-315 4.75121e-315
13425 0
2 5e-005 10
8
199 103
0 12 0 -72 1	0 18 0 0
203 94
0 13 0 -50 1	0 19 0 0
203 85
0 14 0 -29 1	0 20 0 0
206 76
0 15 0 -10 1	0 21 0 0
325 85
0 11 0 16 1	0 17 0 0
330 94
0 10 0 35 1	0 16 0 0
334 112
0 9 0 55 1	0 15 0 0
339 121
0 8 0 71 1	0 14 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
