CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 12 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
70 110 30 200 9
34 91 1332 708
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
53 C:\Users\Josefa Ramos\Documents\Circuit Maker\BOM.DAT
0 7
34 91 1332 708
143654930 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 133 307 0 1 11
0 7
0
0 0 21088 0
2 0V
-6 -16 8 -8
1 D
-3 -17 4 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 133 260 0 1 11
0 11
0
0 0 21088 0
2 0V
-6 -16 8 -8
1 C
-3 -16 4 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 134 219 0 1 11
0 5
0
0 0 21088 0
2 0V
-6 -16 8 -8
1 B
-3 -18 4 -10
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 134 181 0 1 11
0 8
0
0 0 21088 0
2 0V
-6 -16 8 -8
1 A
-4 -17 3 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
14 Logic Display~
6 583 218 0 1 2
12 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 586 347 0 1 2
12 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
9 Inverter~
13 268 338 0 2 22
0 8 6
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
9914 0 0
0
0
9 Inverter~
13 221 213 0 2 22
0 5 13
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3747 0 0
0
0
8 2-In OR~
219 516 365 0 3 22
0 4 7 2
0
0 0 608 0
6 74LS32
-21 -24 21 -16
2 F2
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3549 0 0
0
0
8 2-In OR~
219 516 236 0 3 22
0 10 9 3
0
0 0 608 0
6 74LS32
-21 -24 21 -16
2 F1
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7931 0 0
0
0
9 2-In AND~
219 355 347 0 3 22
0 6 5 4
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9325 0 0
0
0
9 2-In XOR~
219 395 298 0 3 22
0 5 7 9
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 XOR
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8903 0 0
0
0
9 2-In AND~
219 281 222 0 3 22
0 13 11 12
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3834 0 0
0
0
8 2-In OR~
219 389 190 0 3 22
0 8 12 10
0
0 0 608 0
0
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3363 0 0
0
0
16
3 1 2 0 0 4224 0 9 6 0 0 2
549 365
586 365
3 1 3 0 0 4224 0 10 5 0 0 2
549 236
583 236
3 1 4 0 0 4224 0 11 9 0 0 4
376 347
466 347
466 356
503 356
0 2 5 0 0 8192 0 0 11 15 0 3
175 213
175 356
331 356
2 1 6 0 0 4224 0 7 11 0 0 2
289 338
331 338
0 2 7 0 0 8320 0 0 9 10 0 3
217 307
217 374
503 374
0 1 8 0 0 4096 0 0 7 16 0 3
162 181
162 338
253 338
3 2 9 0 0 8320 0 12 10 0 0 4
428 298
460 298
460 245
503 245
3 1 10 0 0 12416 0 14 10 0 0 4
422 190
460 190
460 227
503 227
1 2 7 0 0 0 0 1 12 0 0 2
145 307
379 307
0 1 5 0 0 8320 0 0 12 15 0 3
187 213
187 289
379 289
1 2 11 0 0 4224 0 2 13 0 0 4
145 260
210 260
210 231
257 231
3 2 12 0 0 4224 0 13 14 0 0 4
302 222
339 222
339 199
376 199
2 1 13 0 0 4224 0 8 13 0 0 2
242 213
257 213
1 1 5 0 0 0 0 3 8 0 0 3
146 219
146 213
206 213
1 1 8 0 0 4224 0 4 14 0 0 2
146 181
376 181
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 35
245 134 533 158
250 138 530 154
35 QUEST�O 10 - 2 SA�DAS COM PORTAS OR
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
