CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 640 452
7 5.000 V
7 5.000 V
3 GND
10000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 452
9961472 0
0
0
0
0
0
0
45
2 +V
167 425 306 0 1 64
0 6
0
0 0 54112 0
4 -12V
-15 -14 13 -6
3 Vee
-9 -25 12 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
2 +V
167 150 257 0 1 64
0 7
0
0 0 54112 0
4 +12V
-14 -14 14 -6
3 Vcc
-9 -24 12 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
7 Ground~
168 19 346 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
7 Ground~
168 588 358 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
7 Ground~
168 82 63 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
11 Signal Gen~
195 40 40 0 19 64
0 10 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1036831949 1176256512 0 1036831949
20
0.1 10000 0 0.1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 576 0
11 -100m/100mV
-36 -48 41 -40
3 Vin
-10 -28 11 -20
0
0
43 %D %1 %2 DC 0 SIN(0 100m 10k 0 0) AC 100m 0
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
7 Ground~
168 377 282 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
7 Ground~
168 239 249 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
7 Ground~
168 274 116 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
7 Ground~
168 428 188 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
7 Ground~
168 257 349 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
7 Ground~
168 472 188 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
7 Ground~
168 445 28 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
9 V Source~
197 464 283 0 2 64
0 17 6
0
0 0 17216 0
4 2.6V
12 2 40 10
2 VE
13 -8 27 0
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
2 Vs
3363 0 0
0
0
6 Diode~
219 518 206 0 2 64
0 8 18
6 Diode~
0 0 576 0
5 1N914
-17 -18 18 -10
2 DC
-7 -21 7 -13
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
7668 0 0
0
0
6 Diode~
219 472 110 0 2 64
0 3 4
6 Diode~
0 0 576 270
5 1N914
-17 -18 18 -10
3 DLP
13 -4 34 4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
4718 0 0
0
0
6 Diode~
219 486 321 0 2 64
0 6 7
6 Diode~
0 0 576 0
5 1N914
-17 -18 18 -10
2 DP
-7 -18 7 -10
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
3874 0 0
0
0
6 Diode~
219 481 245 0 2 64
0 17 8
6 Diode~
0 0 576 0
5 1N914
-17 -18 18 -10
2 DE
-7 -20 7 -12
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
6671 0 0
0
0
6 Diode~
219 472 76 0 2 64
0 5 3
6 Diode~
0 0 576 270
5 1N914
-17 -18 18 -10
3 DLN
14 -4 35 4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
3789 0 0
0
0
10 NPN Trans~
219 54 266 0 3 64
0 11 9 14
10 NPN Trans~
0 0 576 0
7 2N2222A
8 -4 57 4
2 Q1
6 -4 20 4
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 -33686019
81 0 0 0 1 1 0 0
1 Q
4871 0 0
0
0
10 NPN Trans~
219 170 302 0 3 64
0 12 2 13
10 NPN Trans~
0 0 576 0
7 2N2222A
8 -4 57 4
2 Q2
5 -4 19 4
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 -33686019
81 0 0 0 1 1 0 0
1 Q
3750 0 0
0
0
9 V Source~
197 472 37 0 2 64
0 2 5
0
0 0 17216 0
3 25V
15 2 36 10
3 VLN
15 -9 36 -1
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
2 Vs
8778 0 0
0
0
9 V Source~
197 472 149 0 2 64
0 4 2
0
0 0 17216 0
3 25V
15 2 36 10
3 VLP
15 -9 36 -1
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
2 Vs
538 0 0
0
0
9 V Source~
197 550 252 0 2 64
0 7 18
0
0 0 17216 180
4 2.6V
12 2 40 10
2 VC
13 -8 27 0
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
2 Vs
6843 0 0
0
0
9 V Source~
197 257 313 0 2 64
0 15 2
0
0 0 17216 0
2 0V
13 4 27 12
2 VB
13 -6 27 2
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
2 Vs
3136 0 0
0
0
12 I->V Source~
201 408 144 0 4 64
0 3 2 21 19
0
0 0 17216 0
2 1K
-8 -19 6 -11
4 HLIM
-12 11 16 19
0
0
32 V%D %3 %4 DC 0V
%D %1 %2 V%D %V
0
0
0
9

0 3 4 1 2 3 4 1 2 -33686019
72 0 0 0 1 0 0 0
4 IcVs
5950 0 0
0
0
9 I Source~
198 312 320 0 2 64
0 16 6
0
0 0 17216 0
8 10.16E-6
11 2 67 10
3 IEE
17 -8 38 0
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 -33686019
73 0 0 0 1 0 0 0
2 Is
5670 0 0
0
0
12 V->I Source~
200 226 120 0 4 64
0 2 22 16 20
0
0 0 17216 0
8 2.574E-9
-20 -19 36 -11
3 GCM
-10 11 11 19
0
0
17 %D %1 %2 %3 %4 %V
0
0
0
9

0 3 4 1 2 3 4 1 2 -33686019
71 0 0 0 1 0 0 0
4 VcIs
6828 0 0
0
0
12 V->I Source~
200 219 207 0 4 64
0 22 2 11 12
0
0 0 17216 0
8 137.7E-6
-20 -19 36 -11
2 GA
-8 11 6 19
0
0
17 %D %1 %2 %3 %4 %V
0
0
0
9

0 3 4 1 2 3 4 1 2 -33686019
71 0 0 0 1 0 0 0
4 VcIs
6735 0 0
0
0
11 NLI Source~
204 331 151 0 2 64
0 21 20
0
0 0 16960 0
5 100mA
-17 -31 18 -23
2 BB
14 -3 28 5
0
0
70 %D %1 %2 I=I(VB)*10.61E6-I(VC)*10E6+I(VE)*10E6+I(VLP)*10E6-I(VLN)*10E6
0
0
0
5

0 1 2 1 2 -33686019
66 0 0 0 1 0 0 0
4 NLIs
8365 0 0
0
0
11 NLV Source~
203 415 247 0 2 64
0 20 2
0
0 0 17216 0
15 V(7)*.5+V(6)*.5
-116 -11 -11 -3
4 BGND
-41 0 -13 8
0
0
13 %D %1 %2 V=%L
0
0
0
5

0 1 2 1 2 -33686019
66 0 0 0 1 0 0 0
4 NLVs
4132 0 0
0
0
10 Polar Cap~
219 80 165 0 2 64
0 11 12
10 Polar Cap~
0 0 832 270
7 4.664pF
10 0 59 8
2 C1
12 -9 26 -1
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
4551 0 0
0
0
10 Polar Cap~
219 278 168 0 2 64
0 22 21
10 Polar Cap~
0 0 832 0
4 20pF
-15 -18 13 -10
2 C2
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3635 0 0
0
0
9 Resistor~
219 484 358 0 3 64
0 6 7 1
9 Resistor~
0 0 4960 0
6 18.11K
-21 -12 21 -4
2 RP
-8 -22 6 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3973 0 0
0
0
9 Resistor~
219 342 96 0 2 64
0 21 20
9 Resistor~
0 0 4960 0
3 150
-11 -12 10 -4
3 RO2
-11 -22 10 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3851 0 0
0
0
9 Resistor~
219 453 219 0 2 64
0 19 8
9 Resistor~
0 0 4960 0
3 150
-11 -12 10 -4
3 RO1
-11 -22 10 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8383 0 0
0
0
9 Resistor~
219 337 225 0 2 64
0 16 20
9 Resistor~
0 0 4960 0
8 19.69Meg
-28 -12 28 -4
3 REE
-11 -22 10 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
9334 0 0
0
0
9 Resistor~
219 127 119 0 2 64
0 13 16
9 Resistor~
0 0 4960 0
5 2.74K
-18 -12 17 -4
3 RE2
-11 -22 10 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7471 0 0
0
0
9 Resistor~
219 128 86 0 2 64
0 14 16
9 Resistor~
0 0 4960 0
5 2.74K
-18 -12 17 -4
3 RE1
-11 -22 10 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3334 0 0
0
0
9 Resistor~
219 127 208 0 3 64
0 7 12 1
9 Resistor~
0 0 4960 90
6 7.957K
5 3 47 11
3 RC2
6 -9 27 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3559 0 0
0
0
9 Resistor~
219 257 264 0 2 64
0 15 22
9 Resistor~
0 0 4960 90
4 100k
5 4 33 12
2 R2
7 -6 21 2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
984 0 0
0
0
9 Resistor~
219 94 236 0 4 64
0 11 7 0 1
9 Resistor~
0 0 4960 0
6 7.957K
-21 -12 21 -4
3 RC1
-11 -22 10 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7557 0 0
0
0
9 Resistor~
219 118 35 0 2 64
0 10 9
9 Resistor~
0 0 4960 0
3 10k
-10 -12 11 -4
2 RI
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3146 0 0
0
0
9 Resistor~
219 196 35 0 2 64
0 9 8
9 Resistor~
0 0 4960 0
4 100k
-14 -12 14 -4
2 RF
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
5687 0 0
0
0
9 Resistor~
219 559 345 0 4 64
0 8 2 0 -1
9 Resistor~
0 0 4960 0
3 25k
-10 -12 11 -4
2 RL
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7939 0 0
0
0
56
1 0 3 0 0 8320 0 26 0 0 3 3
428 117
428 93
472 93
2 1 4 0 0 12416 0 16 23 0 0 4
472 120
472 119
472 119
472 128
2 1 3 0 0 0 0 19 16 0 0 2
472 86
472 100
2 1 5 0 0 4224 0 22 19 0 0 2
472 58
472 66
1 0 6 0 0 4096 0 1 0 0 30 2
425 315
425 348
1 0 7 0 0 8192 0 2 0 0 28 3
150 266
150 276
127 276
2 0 8 0 0 16512 0 44 0 0 8 6
214 35
312 35
312 7
602 7
602 315
533 315
0 1 8 0 0 0 0 0 45 37 0 4
498 233
533 233
533 345
541 345
2 1 2 0 0 4096 0 45 4 0 0 3
577 345
588 345
588 352
0 2 9 0 0 12416 0 0 20 11 0 5
150 35
150 6
8 6
8 266
48 266
2 1 9 0 0 0 0 43 44 0 0 2
136 35
178 35
1 1 10 0 0 4224 0 6 43 0 0 2
71 35
100 35
2 1 2 0 0 8192 0 6 5 0 0 3
71 45
82 45
82 57
2 1 2 0 0 4224 0 21 3 0 0 3
164 302
19 302
19 340
1 0 11 0 0 4096 0 32 0 0 56 2
79 155
79 146
2 0 7 0 0 0 0 42 0 0 28 2
112 236
127 236
2 0 12 0 0 4096 0 40 0 0 54 2
127 190
127 179
1 1 2 0 0 0 0 28 9 0 0 3
246 93
274 93
274 110
2 1 2 0 0 0 0 26 10 0 0 2
428 171
428 182
2 1 2 0 0 0 0 29 8 0 0 2
239 234
239 243
1 1 2 0 0 0 0 22 13 0 0 4
472 16
472 10
445 10
445 22
2 1 2 0 0 0 0 23 12 0 0 2
472 170
472 182
2 1 2 0 0 0 0 31 7 0 0 4
415 268
415 272
377 272
377 276
2 1 2 0 0 0 0 25 11 0 0 2
257 334
257 343
3 1 13 0 0 12416 0 21 38 0 0 5
177 320
177 333
29 333
29 119
109 119
3 1 14 0 0 12416 0 20 39 0 0 5
61 284
61 291
38 291
38 86
110 86
0 1 7 0 0 8192 0 0 24 32 0 4
515 321
515 302
550 302
550 271
0 1 7 0 0 8320 0 0 40 32 0 4
515 357
515 368
127 368
127 226
1 1 15 0 0 4224 0 41 25 0 0 2
257 282
257 292
2 0 6 0 0 8320 0 27 0 0 33 3
312 341
312 348
449 348
0 1 16 0 0 4096 0 0 27 41 0 4
293 225
293 284
312 284
312 299
2 2 7 0 0 0 0 17 34 0 0 4
496 321
515 321
515 358
502 358
0 1 6 0 0 0 0 0 34 34 0 4
464 321
449 321
449 358
466 358
2 1 6 0 0 0 0 14 17 0 0 3
464 304
464 321
476 321
1 1 17 0 0 8320 0 18 14 0 0 3
471 245
464 245
464 262
2 2 18 0 0 4224 0 24 15 0 0 3
550 229
550 206
528 206
2 0 8 0 0 0 0 18 0 0 38 3
491 245
498 245
498 219
2 1 8 0 0 0 0 36 15 0 0 4
471 219
498 219
498 206
508 206
4 1 19 0 0 4224 0 26 36 0 0 3
388 171
388 219
435 219
2 1 20 0 0 8192 0 30 31 0 0 4
331 172
331 184
415 184
415 226
0 1 16 0 0 8320 0 0 37 43 0 4
206 86
293 86
293 225
319 225
2 0 16 0 0 0 0 38 0 0 43 3
145 119
163 119
163 86
2 3 16 0 0 0 0 39 28 0 0 3
146 86
206 86
206 93
0 4 20 0 0 8320 0 0 28 45 0 6
368 96
368 67
177 67
177 153
206 153
206 147
2 0 20 0 0 0 0 35 0 0 46 3
360 96
368 96
368 184
2 0 20 0 0 0 0 37 0 0 40 3
355 225
368 225
368 184
0 3 21 0 0 4224 0 0 26 49 0 3
331 112
388 112
388 117
1 0 21 0 0 0 0 35 0 0 49 3
324 96
317 96
317 112
2 1 21 0 0 0 0 33 30 0 0 5
284 168
306 168
306 112
331 112
331 130
2 0 22 0 0 4224 0 41 0 0 52 2
257 246
257 168
2 0 22 0 0 0 0 28 0 0 52 2
246 147
246 168
1 1 22 0 0 0 0 33 29 0 0 3
267 168
239 168
239 180
4 0 12 0 0 8192 0 29 0 0 54 3
199 234
199 240
177 240
2 1 12 0 0 12416 0 32 21 0 0 4
79 172
79 179
177 179
177 284
0 1 11 0 0 4096 0 0 42 56 0 2
61 236
76 236
3 1 11 0 0 20608 0 29 20 0 0 6
199 180
199 168
160 168
160 146
61 146
61 248
0
0
17 0 0
0
0
3 Vin
-1.5 -0.7 0.01
3 Vcc
10 14 1
100 0 1 100000
0 0.0005 2.5e-006 2.5e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
