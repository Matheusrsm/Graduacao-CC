CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 100 9
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
5000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 259
9961474 0
0
0
0
0
0
0
3
7 Ground~
168 165 173 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
11 Signal Gen~
195 87 141 0 32 64
0 3 2 5 86 -8 8 9 0 0
0 0 0 0 0 0 0 0 0 0
897988541 0 906377149 1065353216 910775196 1073741824 914765757 -1090519040 916964780 1056964608
919163804 0 921362827
20
0 0 0 0 1e-006 0 2e-006 1 3e-006 2
4e-006 -0.5 5e-006 0.5 6e-006 0 7e-006 0 0 0
0
0 0 832 0
4 0/0V
-14 -28 14 -20
2 V1
-7 -38 7 -30
0
0
44 %D %1 %2 DC 0 PWL %=RAND128.PWL{0.5 0.001 1}
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
9 Resistor~
219 186 121 0 4 64
0 3 2 0 -1
9 Resistor~
0 0 864 0
2 1k
-7 -12 7 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3618 0 0
0
0
3
1 0 2 0 0 4096 0 1 0 0 2 2
165 167
165 154
2 2 2 0 0 12416 0 2 3 0 0 6
118 146
131 146
131 154
234 154
234 121
204 121
1 1 3 0 0 4224 0 3 2 0 0 4
168 121
131 121
131 136
118 136
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 152
7 38 430 102
11 42 427 94
152 This circuit demonstrates the use of a piece-wise 
linear signal generator whose output is determined 
from an external data file named RAND128.PWL.
0
16 0 1
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 0.001 2.5e-005 2.5e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3272 8550464 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 67
617 126
0 0
4.85009e-315 0 5.271e-315 0 4.85009e-315 4.85009e-315
0 0
4 0.0002 0.5
1
152 121
0 3 0 0 1	0 3 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
