CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 640 452
7 5.000 V
7 5.000 V
3 GND
0 66 640 452
9437184 0
0
0
0
0
0
0
18
9 Inverter~
13 359 231 0 2 21
0 26 4
0
0 0 112 90
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 2 1 0
1 U
8953 0 0
0
0
14 Logic Display~
6 293 33 0 1 3
10 6
0
0 0 53344 0
6 100MEG
3 -16 45 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
13 Piezo Buzzer~
174 480 223 0 2 5
10 5 2
0
0 0 4208 270
4 .1uF
10 -16 38 -8
0
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
2 BZ
3618 0 0
0
0
8 Hex Key~
166 362 45 0 11 11
0 9 10 11 12 0 0 0 0 0
0 48
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6153 0 0
0
0
8 Hex Key~
166 326 45 0 11 11
0 13 14 15 16 0 0 0 0 0
8 56
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5394 0 0
0
0
5 Delay
94 416 104 0 11 23
0 16 15 14 13 12 11 10 9 5
8 7
5 Delay
1 0 4240 0
0
0
0
0
0
0
0
0
23

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
7 Ground~
168 232 282 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
8 Hex Key~
166 76 44 0 11 11
0 18 19 20 21 0 0 0 0 0
0 48
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3747 0 0
0
0
8 Hex Key~
166 38 44 0 11 11
0 22 23 24 25 0 0 0 0 0
4 52
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3549 0 0
0
0
5 Delay
94 129 105 0 11 23
0 25 24 23 22 21 20 19 18 6
17 7
5 Delay
2 0 4240 0
0
0
0
0
0
0
0
0
23

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
6 74LS74
17 417 214 0 12 25
0 85 86 4 6 87 88 89 90 91
8 92 93
0
0 0 12464 0
6 74LS74
-21 -60 21 -52
0
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 -33686019
65 0 0 512 1 1 0 0
1 U
9325 0 0
0
0
14 NO PushButton~
191 259 124 0 2 5
0 17 2
0
0 0 20592 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8903 0 0
0
0
14 NO PushButton~
191 207 124 0 2 5
0 2 7
0
0 0 20592 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3834 0 0
0
0
7 Window~
179 270 217 0 4 9
0 26 6 94 95
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 WND
3363 0 0
0
0
7 Ground~
168 480 278 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
7 Window~
179 146 217 0 4 9
0 26 6 96 97
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 WND
4718 0 0
0
0
7 Window~
179 37 218 0 4 9
0 26 6 98 99
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 WND
3874 0 0
0
0
9 Resistor~
219 406 265 0 4 64
0 26 2 0 -1
9 Resistor~
0 0 4208 0
2 1k
-7 -14 7 -6
0
0
0
11 %D %1 %2 %V
0
0
0
3

0 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
35
1 0 2 0 0 4224 0 7 0 0 18 2
232 276
232 132
2 3 4 0 0 4224 0 1 11 0 0 3
362 213
362 196
379 196
2 0 2 0 0 0 0 18 0 0 5 2
424 265
480 265
1 9 5 0 0 4224 0 3 6 0 0 3
480 192
480 86
448 86
2 1 2 0 0 0 0 3 15 0 0 2
480 254
480 272
1 0 6 0 0 4096 0 2 0 0 23 2
293 51
293 163
0 11 7 0 0 8320 0 0 6 20 0 5
180 132
180 155
468 155
468 131
454 131
10 10 8 0 0 8320 0 6 11 0 0 4
454 140
461 140
461 196
455 196
8 1 9 0 0 8320 0 6 4 0 0 3
384 140
371 140
371 69
2 7 10 0 0 4224 0 4 6 0 0 3
365 69
365 131
384 131
3 6 11 0 0 4224 0 4 6 0 0 3
359 69
359 122
384 122
5 4 12 0 0 8320 0 6 4 0 0 3
384 113
353 113
353 69
1 4 13 0 0 8320 0 5 6 0 0 3
335 69
335 104
384 104
2 3 14 0 0 8320 0 5 6 0 0 3
329 69
329 95
384 95
3 2 15 0 0 8320 0 5 6 0 0 3
323 69
323 86
384 86
1 4 16 0 0 4224 0 6 5 0 0 3
384 77
317 77
317 69
4 0 6 0 0 0 0 11 0 0 23 2
379 205
325 205
2 1 2 0 0 0 0 12 13 0 0 2
242 132
224 132
10 1 17 0 0 4224 0 10 12 0 0 4
167 141
287 141
287 132
276 132
11 2 7 0 0 0 0 10 13 0 0 2
167 132
190 132
9 0 6 0 0 0 0 10 0 0 23 3
161 87
172 87
172 163
2 0 6 0 0 0 0 16 0 0 23 3
192 226
205 226
205 163
2 2 6 0 0 12416 0 14 17 0 0 6
316 226
325 226
325 163
94 163
94 227
83 227
8 1 18 0 0 8320 0 10 8 0 0 3
97 141
85 141
85 68
2 7 19 0 0 4224 0 8 10 0 0 3
79 68
79 132
97 132
3 6 20 0 0 4224 0 8 10 0 0 3
73 68
73 123
97 123
5 4 21 0 0 8320 0 10 8 0 0 3
97 114
67 114
67 68
1 4 22 0 0 8320 0 9 10 0 0 3
47 68
47 105
97 105
2 3 23 0 0 8320 0 9 10 0 0 3
41 68
41 96
97 96
3 2 24 0 0 8320 0 9 10 0 0 3
35 68
35 87
97 87
1 4 25 0 0 4224 0 10 9 0 0 3
97 78
29 78
29 68
1 1 26 0 0 12416 0 17 18 0 0 4
83 236
95 236
95 265
388 265
1 0 26 0 0 0 0 16 0 0 32 3
192 235
205 235
205 265
1 0 26 0 0 0 0 1 0 0 32 2
362 249
362 265
1 0 26 0 0 0 0 14 0 0 32 3
316 235
326 235
326 265
5
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 5
229 22 288 49
233 26 278 45
5 Armed
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 13
231 67 298 117
235 71 288 109
13 Enable
Alarm
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 12
179 67 246 117
183 71 236 109
12 Reset
Alarm
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 16
97 18 182 68
101 22 172 60
16 Exit Delay
Time
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 19
389 18 488 68
393 22 478 60
19 Entry Delay 
Time
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 100 100 0 0
77 66 617 126
0 0 0 0
617 66
77 66
617 66
617 126
0 0
0.0005 0 1.2 -1.2 0.0005 0.0005
16 0
0 0.0001 10
0
0 0 100 100 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 -1.#IND -1.#IND 0 0
0 0
0 0.0002 10
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
