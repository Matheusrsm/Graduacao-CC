CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 12 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
210 80 30 200 9
93 93 1333 746
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 Z:\home\matheussm\Documentos\UFCG\P1\IC\Circuit Maker\BOM.DAT
0 7
93 93 1333 746
143654930 0
0
6 Title:
5 Name:
0
0
0
7
13 Logic Switch~
5 327 297 0 1 11
0 2
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 A
-4 -17 3 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 327 248 0 1 11
0 6
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 C
-3 -16 4 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 326 206 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
1 B
-3 -16 4 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
14 Logic Display~
6 616 228 0 1 2
12 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
9 Inverter~
13 451 204 0 2 22
0 8 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
5394 0 0
0
0
9 2-In AND~
219 439 275 0 3 22
0 6 3 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7734 0 0
0
0
8 2-In OR~
219 549 246 0 3 22
0 7 5 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
2 OR
-1 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9914 0 0
0
0
6
1 2 3 0 0 8336 0 1 6 0 0 3
339 297
339 284
415 284
3 1 4 0 0 4224 0 7 4 0 0 2
582 246
616 246
3 2 5 0 0 4224 0 6 7 0 0 4
460 275
510 275
510 255
536 255
1 1 6 0 0 8320 0 2 6 0 0 3
339 248
339 266
415 266
2 1 7 0 0 8320 0 5 7 0 0 3
472 204
472 237
536 237
1 1 8 0 0 8320 0 3 5 0 0 3
338 206
338 204
436 204
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 38
401 137 562 181
405 139 558 171
38  QUEST�O 6(ITEM B)
SA�DA COM PORTA OR
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
