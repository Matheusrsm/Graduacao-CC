CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 90 9 100 9
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
1.66667 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 259
11010066 0
0
0
0
0
0
0
15
11 Signal Gen~
195 38 133 0 64 64
0 3 2 1 86 -8 8 0 0 0
0 0 0 0 0 0 0 1065353216 0 1083179008
1056964608 1020054733 1020054733 1045220557 1065353216 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
20
0 1 0 4.5 0.5 0.025 0.025 0.2 1 0
0 0 0 0 0 0 0 0 0 0
0
0 0 320 0
6 0/4.5V
-20 -28 22 -20
2 V1
-7 -38 7 -30
0
0
46 %D %1 %2 DC 0 PULSE(0 4.5 500m 25m 25m 200m 1)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
9 2-In NOR~
219 383 173 0 3 21
0 5 5 4
0
0 0 96 0
6 74LS02
-21 -24 21 -16
3 U1B
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 2 1 0
1 U
4441 0 0
0
0
9 2-In NOR~
219 290 164 0 3 21
0 7 6 5
0
0 0 96 0
6 74LS02
-21 -24 21 -16
3 U1A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 1 0
1 U
3618 0 0
0
0
4 .IC~
207 234 175 0 1 3
0 6
0
0 0 53568 0
2 0V
-7 -15 7 -7
4 CMD1
-14 -25 14 -17
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
3 CMD
6153 0 0
0
0
12 SPST Switch~
165 327 192 0 2 11
0 6 4
0
0 0 20576 512
0
2 S1
-7 -28 7 -20
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5394 0 0
0
0
7 Ground~
168 77 150 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
2 +V
167 207 96 0 1 3
0 8
0
0 0 53600 0
3 +5V
12 -2 33 6
2 V2
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
7 Ground~
168 194 244 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
4 LED~
171 482 211 0 2 5
12 5 9
0
0 0 608 0
4 LED2
10 -16 38 -8
2 D1
17 -26 31 -18
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3549 0 0
0
0
4 LED~
171 431 211 0 2 5
10 4 9
0
0 0 608 0
4 LED2
10 -16 38 -8
2 D2
17 -26 31 -18
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7931 0 0
0
0
12 NPN Trans:C~
219 202 128 0 3 7
0 8 10 7
12 NPN Trans:C~
0 0 832 0
6 2N3904
20 -4 62 4
2 Q1
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
9325 0 0
0
0
9 Resistor~
219 388 237 0 3 11
0 2 9 -1
9 Resistor~
0 0 864 0
3 150
-10 -12 11 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 256 216 0 3 11
0 2 6 -1
9 Resistor~
0 0 864 90
3 470
4 3 25 11
2 R2
6 -7 20 1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 207 212 0 3 11
0 2 7 -1
9 Resistor~
0 0 864 90
3 470
7 1 28 9
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 152 128 0 2 11
0 3 10
9 Resistor~
0 0 864 0
2 1k
-7 -12 7 -4
2 R4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
7668 0 0
0
0
19
2 1 2 0 0 4096 0 1 6 0 0 3
69 138
77 138
77 144
1 1 3 0 0 4224 0 15 1 0 0 2
134 128
69 128
3 1 4 0 0 8192 0 2 10 0 0 3
422 173
431 173
431 201
1 2 5 0 0 4096 0 2 2 0 0 4
370 164
349 164
349 182
370 182
3 0 5 0 0 0 0 3 0 0 4 2
329 164
349 164
2 2 6 0 0 8192 0 3 13 0 0 3
277 173
256 173
256 198
1 0 7 0 0 4224 0 3 0 0 18 2
277 155
207 155
1 0 2 0 0 8192 0 8 0 0 17 3
194 238
194 237
207 237
1 0 6 0 0 0 0 4 0 0 6 3
234 187
234 192
256 192
1 0 5 0 0 8320 0 9 0 0 5 4
482 201
482 127
349 127
349 164
1 0 6 0 0 4224 0 5 0 0 6 2
310 192
256 192
2 0 4 0 0 4224 0 5 0 0 3 2
344 192
431 192
1 1 8 0 0 4224 0 7 11 0 0 2
207 105
207 110
2 0 9 0 0 4096 0 10 0 0 15 2
431 221
431 237
2 2 9 0 0 4224 0 12 9 0 0 3
406 237
482 237
482 221
1 0 2 0 0 0 0 13 0 0 17 2
256 234
256 237
1 1 2 0 0 8320 0 14 12 0 0 3
207 230
207 237
370 237
3 2 7 0 0 0 0 11 14 0 0 2
207 146
207 194
2 2 10 0 0 4224 0 15 11 0 0 2
170 128
184 128
2
-11 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
97 129 167 149
101 133 164 147
9 Probe Tip
-20 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 11
347 90 488 125
351 94 483 121
11 Logic Probe
19 .OPTIONS TRTOL=10

16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 3 0.025 0.025
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
164 8526400 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 89
617 98
0 0
5.32571e-315 0 5.33607e-315 1.58735e-314 5.32571e-315 5.32571e-315
13433 0
2 0.5 5
3
109 128
0 3 0 16 1	0 2 0 0
482 168
0 5 0 0 1	0 10 0 0
431 173
0 4 0 -15 1	0 3 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
