CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 200 9
63 134 1370 772
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
54 C:\Users\H�rcules\Desktop\Circuito Maker\CM60S\BOM.DAT
0 7
63 134 1370 772
210763794 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 218 36 0 1 11
0 9
0
0 0 21344 0
2 0V
-5 -16 9 -8
2 D2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 348 45 0 1 11
0 11
0
0 0 21344 0
2 0V
-5 -16 9 -8
2 D1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 82 42 0 1 11
0 13
0
0 0 21344 0
2 0V
-5 -16 9 -8
2 D3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 480 51 0 1 11
0 15
0
0 0 21344 0
2 0V
-5 -16 9 -8
2 D0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 53 172 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
5 CLOCK
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 50 222 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
5 CLEAR
-17 -26 18 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7734 0 0
0
0
6 JK RN~
219 286 92 0 6 22
0 9 6 8 5 16 4
0
0 0 4192 0
6 74LS73
-22 -42 20 -34
3 U5A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 10 0
1 U
9914 0 0
0
0
9 Inverter~
13 236 72 0 2 22
0 9 8
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 no2A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 9 0
1 U
3747 0 0
0
0
6 JK RN~
219 416 101 0 6 22
0 11 6 10 5 17 3
0
0 0 4192 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 8 0
1 U
3549 0 0
0
0
9 Inverter~
13 366 81 0 2 22
0 11 10
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 no1F
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 6 6 0
1 U
7931 0 0
0
0
14 Logic Display~
6 449 44 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 183 44 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 325 42 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
0
0
9 Inverter~
13 100 78 0 2 22
0 13 12
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 no1D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 6 0
1 U
3363 0 0
0
0
6 JK RN~
219 150 98 0 6 22
0 13 6 12 5 18 7
0
0 0 4192 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 7 0
1 U
7668 0 0
0
0
14 Logic Display~
6 604 47 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
9 Inverter~
13 499 91 0 2 22
0 15 14
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 no1A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 6 0
1 U
3874 0 0
0
0
6 JK RN~
219 568 119 0 6 22
0 15 6 14 5 19 2
0
0 0 4192 0
6 74LS73
-22 -42 20 -34
3 U4A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 5 0
1 U
6671 0 0
0
0
25
6 1 2 0 0 8320 0 18 16 0 0 3
592 102
604 102
604 65
6 1 3 0 0 8320 0 9 11 0 0 3
440 84
449 84
449 62
1 6 4 0 0 4224 0 13 7 0 0 3
325 60
325 75
310 75
4 0 5 0 0 4096 0 15 0 0 25 2
150 129
150 222
2 0 6 0 0 4096 0 15 0 0 20 2
119 90
119 173
2 0 6 0 0 4096 0 7 0 0 20 2
255 84
255 173
2 0 6 0 0 0 0 9 0 0 20 2
385 93
385 173
4 0 5 0 0 0 0 9 0 0 25 2
416 132
416 222
4 0 5 0 0 4096 0 7 0 0 25 2
286 123
286 222
1 6 7 0 0 4224 0 12 15 0 0 3
183 62
183 81
174 81
3 2 8 0 0 4224 0 7 8 0 0 4
262 93
238 93
238 90
239 90
1 1 9 0 0 4112 0 8 1 0 0 3
239 54
239 36
230 36
1 1 9 0 0 4224 0 8 7 0 0 3
239 54
262 54
262 75
3 2 10 0 0 4224 0 9 10 0 0 4
392 102
368 102
368 99
369 99
1 1 11 0 0 4096 0 10 2 0 0 3
369 63
369 45
360 45
1 1 11 0 0 4224 0 10 9 0 0 3
369 63
392 63
392 84
3 2 12 0 0 4224 0 15 14 0 0 4
126 99
102 99
102 96
103 96
1 1 13 0 0 4096 0 14 3 0 0 3
103 60
103 42
94 42
1 1 13 0 0 4224 0 14 15 0 0 3
103 60
126 60
126 81
0 1 6 0 0 4224 0 0 5 0 0 3
531 173
65 173
65 172
2 0 6 0 0 0 0 18 0 0 20 3
537 111
528 111
528 173
3 2 14 0 0 4224 0 18 17 0 0 3
544 120
502 120
502 109
1 1 15 0 0 4096 0 17 4 0 0 3
502 73
502 51
492 51
1 1 15 0 0 4224 0 17 18 0 0 3
502 73
544 73
544 102
1 4 5 0 0 4224 0 6 18 0 0 3
62 222
568 222
568 150
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
