CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 20 9 100 9
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
5e+006 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 259
11010054 0
0
0
0
0
0
0
27
13 Logic Switch~
5 87 222 0 1 11
0 18
0
0 0 4448 0
2 0V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 87 194 0 1 11
0 19
0
0 0 4448 0
2 0V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
9 Inverter~
13 549 316 0 2 21
0 6 12
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 2 8 0
1 U
3618 0 0
0
0
9 Inverter~
13 547 268 0 2 21
0 7 11
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 1 8 0
1 U
6153 0 0
0
0
9 Inverter~
13 547 223 0 2 21
0 13 10
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U2F
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 6 5 0
1 U
5394 0 0
0
0
9 Inverter~
13 546 178 0 2 21
0 3 9
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 5 5 0
1 U
7734 0 0
0
0
10 2-In NAND~
219 141 203 0 3 21
0 19 18 8
0
0 0 96 0
6 74LS00
-14 -24 28 -16
3 U4A
-4 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 7 0
1 U
9914 0 0
0
0
6 74112~
219 460 152 0 7 31
0 5 5 7 5 8 21 6
0
0 0 4192 0
7 74LS112
-3 -60 46 -52
3 U3B
11 -70 32 -62
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -33686019
65 0 0 512 2 2 6 0
1 U
3747 0 0
0
0
6 74112~
219 365 152 0 7 31
0 5 5 13 5 8 22 7
0
0 0 4192 0
7 74LS112
-3 -60 46 -52
3 U3A
11 -70 32 -62
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -33686019
65 0 0 512 2 1 6 0
1 U
3549 0 0
0
0
6 74112~
219 268 151 0 7 31
0 5 5 3 5 8 23 13
0
0 0 4192 0
7 74LS112
-3 -60 46 -52
3 U1B
11 -70 32 -62
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -33686019
65 0 0 512 2 2 4 0
1 U
7931 0 0
0
0
6 74112~
219 178 150 0 7 31
0 5 5 20 5 8 24 3
0
0 0 4192 0
7 74LS112
-3 -60 46 -52
3 U1A
11 -70 32 -62
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -33686019
65 0 0 512 2 1 4 0
1 U
9325 0 0
0
0
2 +V
167 687 63 0 1 3
0 4
0
0 0 53600 0
4 +15V
-14 -14 14 -6
2 V3
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
7 Ground~
168 760 348 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
7 Ground~
168 711 303 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
7 Ground~
168 659 254 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
7 Ground~
168 606 211 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4718 0 0
0
0
2 +V
167 268 56 0 1 3
0 5
0
0 0 53600 0
3 +5V
12 -2 33 6
2 V4
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3874 0 0
0
0
7 Ground~
168 81 153 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
11 Signal Gen~
195 38 128 0 24 64
0 20 2 1 86 -9 9 0 0 0
0 0 0 0 0 0 0 1259902592 0 1084227584
841731191 833342583 833342583 861323157 869711765
20
0 1e+007 0 5 1e-008 5e-009 5e-009 5e-008 1e-007 0
0 0 0 0 0 0 0 0 0 0
0
0 0 320 0
4 0/5V
-14 -28 14 -20
2 V5
-7 -38 7 -30
0
0
43 %D %1 %2 DC 0 PULSE(0 5 10n 5n 5n 50n 100n)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3789 0 0
0
0
12 NPN Trans:C~
219 601 178 0 3 7
0 17 9 2
12 NPN Trans:C~
0 0 320 0
3 NPN
17 -5 38 3
2 Q1
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
4871 0 0
0
0
12 NPN Trans:C~
219 654 223 0 3 7
0 16 10 2
12 NPN Trans:C~
0 0 320 0
3 NPN
17 -5 38 3
2 Q2
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
3750 0 0
0
0
12 NPN Trans:C~
219 706 268 0 3 7
0 15 11 2
12 NPN Trans:C~
0 0 320 0
3 NPN
17 -5 38 3
2 Q3
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
8778 0 0
0
0
12 NPN Trans:C~
219 755 316 0 3 7
0 14 12 2
12 NPN Trans:C~
0 0 320 0
3 NPN
17 -5 38 3
2 Q4
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
538 0 0
0
0
9 Resistor~
219 606 123 0 4 5
0 17 4 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 659 128 0 4 5
0 16 4 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3136 0 0
0
0
9 Resistor~
219 711 130 0 4 5
0 15 4 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
5950 0 0
0
0
9 Resistor~
219 760 131 0 4 5
0 14 4 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
5670 0 0
0
0
43
3 0 3 0 0 4096 0 10 0 0 2 2
238 124
220 124
7 1 3 0 0 12416 0 11 6 0 0 4
202 114
220 114
220 178
531 178
1 0 4 0 0 4096 0 12 0 0 32 2
687 72
687 93
1 0 5 0 0 4096 0 10 0 0 17 2
268 88
268 76
7 1 6 0 0 8320 0 8 3 0 0 4
484 116
501 116
501 316
534 316
0 1 7 0 0 4224 0 0 4 18 0 3
411 125
411 268
532 268
1 0 5 0 0 8192 0 8 0 0 17 3
460 89
460 76
422 76
1 0 5 0 0 0 0 9 0 0 17 2
365 89
365 76
1 0 5 0 0 0 0 11 0 0 17 2
178 87
178 76
1 0 5 0 0 0 0 17 0 0 17 2
268 65
268 76
2 0 5 0 0 0 0 8 0 0 17 2
436 116
422 116
2 0 5 0 0 0 0 9 0 0 13 2
341 116
327 116
4 0 5 0 0 8192 0 9 0 0 17 3
341 134
327 134
327 76
2 0 5 0 0 0 0 10 0 0 15 2
244 115
231 115
4 0 5 0 0 0 0 10 0 0 17 3
244 133
231 133
231 76
2 0 5 0 0 0 0 11 0 0 17 2
154 114
144 114
4 4 5 0 0 12416 0 11 8 0 0 6
154 132
144 132
144 76
422 76
422 134
436 134
7 3 7 0 0 0 0 9 8 0 0 4
389 116
411 116
411 125
430 125
5 0 8 0 0 4096 0 9 0 0 43 2
365 164
365 203
5 0 8 0 0 4096 0 10 0 0 43 2
268 163
268 203
2 2 9 0 0 4224 0 20 6 0 0 2
583 178
567 178
2 2 10 0 0 4224 0 5 21 0 0 2
568 223
636 223
2 2 11 0 0 4224 0 22 4 0 0 2
688 268
568 268
2 2 12 0 0 4224 0 3 23 0 0 2
570 316
737 316
1 0 13 0 0 4224 0 5 0 0 41 3
532 223
315 223
315 125
3 1 2 0 0 4096 0 23 13 0 0 2
760 334
760 342
3 1 2 0 0 4096 0 22 14 0 0 2
711 286
711 297
3 1 2 0 0 0 0 21 15 0 0 2
659 241
659 248
3 1 2 0 0 0 0 20 16 0 0 2
606 196
606 205
2 0 4 0 0 0 0 26 0 0 32 2
711 112
711 93
2 0 4 0 0 0 0 25 0 0 32 2
659 110
659 93
2 2 4 0 0 8320 0 24 27 0 0 4
606 105
606 93
760 93
760 113
1 1 14 0 0 4224 0 27 23 0 0 2
760 149
760 298
1 1 15 0 0 4224 0 26 22 0 0 2
711 148
711 250
1 1 16 0 0 4224 0 25 21 0 0 2
659 146
659 205
1 1 17 0 0 4224 0 24 20 0 0 2
606 141
606 160
1 2 18 0 0 12416 0 1 7 0 0 4
99 222
103 222
103 212
117 212
1 1 19 0 0 4224 0 2 7 0 0 2
99 194
117 194
1 3 20 0 0 4224 0 19 11 0 0 2
69 123
148 123
2 1 2 0 0 8320 0 19 18 0 0 3
69 133
81 133
81 147
7 3 13 0 0 0 0 10 9 0 0 4
292 115
315 115
315 125
335 125
5 0 8 0 0 4096 0 11 0 0 43 2
178 162
178 203
3 5 8 0 0 4224 0 7 8 0 0 3
168 203
460 203
460 164
5
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
502 295 526 319
506 299 522 315
2 Q3
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
500 157 525 181
504 161 520 177
2 Q0
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
500 202 524 226
504 206 520 222
2 Q1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
501 247 526 271
505 251 521 267
2 Q2
-20 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 40
25 16 514 51
29 20 509 47
40 Mixed-mode Binary Ripple Counter Circuit
0
16 0 1
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 1e-006 2.5e-008 2.5e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2744 8522304 100 100 0 0
98 66 608 126
0 259 640 452
606 66
98 66
608 69
608 74
0 0
0 0 0 0 0 0
12409 0
4 3e-007 2
1
108 123
0 20 0 0 1	0 39 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
