CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
16 74 624 456
7 5.000 V
7 5.000 V
3 GND
16 74 624 456
142606338 0
0
0
0
0
0
0
2
13 Logic Switch~
5 105 96 0 2 3
0 2 -99
0
0 0 20576 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 0 0 0 0
1 V
8953 0 0
0
0
9 Inverter~
13 219 96 0 2 21
0 3 4
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 512 6 1 1 0
1 U
4441 0 0
0
0
0
3
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 12
69 106 145 127
73 110 142 125
12 Logic Switch
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 8
196 105 248 129
200 109 249 129
8 Inverter
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 29
117 36 281 57
121 40 278 55
29 Place a Logic Display here =>
0
29 0 1
0
0
3 Vin
-1.5 -0.7 0.01
3 Vcc
10 14 1
100 0 1 1e+006
0 0.0005 2.5e-006 2.5e-006 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
