CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 12 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
300 90 30 400 9
34 91 1332 708
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
53 C:\Users\Josefa Ramos\Documents\Circuit Maker\BOM.DAT
0 7
34 91 1332 708
143654930 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 394 225 0 1 11
0 4
0
0 0 21104 0
2 0V
-6 -16 8 -8
2 T2
-6 -17 8 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 394 186 0 1 11
0 5
0
0 0 21104 0
2 0V
-6 -16 8 -8
2 T1
-6 -18 8 -10
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
14 Logic Display~
6 578 231 0 1 2
12 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 576 162 0 1 2
12 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
9 Inverter~
13 457 194 0 2 22
0 4 6
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
5394 0 0
0
0
9 Inverter~
13 457 166 0 2 22
0 5 7
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
7734 0 0
0
0
9 2-In AND~
219 534 249 0 3 22
0 5 4 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
1 R
-5 -25 2 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9914 0 0
0
0
9 2-In AND~
219 533 180 0 3 22
0 7 6 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
1 A
-5 -25 2 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3747 0 0
0
0
8
3 1 2 0 0 4224 0 7 3 0 0 2
555 249
578 249
3 1 3 0 0 4224 0 8 4 0 0 2
554 180
576 180
0 2 4 0 0 8336 0 0 7 5 0 3
427 225
427 258
510 258
0 1 5 0 0 8320 0 0 7 6 0 3
418 186
418 240
510 240
1 1 4 0 0 0 0 1 5 0 0 4
406 225
436 225
436 194
442 194
1 1 5 0 0 0 0 2 6 0 0 4
406 186
428 186
428 166
442 166
2 2 6 0 0 4224 0 5 8 0 0 4
478 194
501 194
501 189
509 189
2 1 7 0 0 4224 0 6 8 0 0 4
478 166
501 166
501 171
509 171
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 47
390 103 582 147
393 105 577 137
47  COMPLEMENTAR - ESTUFA
2 SA�DAS COM PORTAS AND
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
