logic [6:0] entrada;

always_comb begin
	entrada <= SWI[6:0];
	case(entrada)

		// Números Hexadecimais

		0: SEG[6:0] <= 7'b0111111;
		1: SEG[6:0] <= 7'b0000110;
		2: SEG[6:0] <= 7'b1011011;
		3: SEG[6:0] <= 7'b1001111;
		4: SEG[6:0] <= 7'b1100110;
		5: SEG[6:0] <= 7'b1101101;
		6: SEG[6:0] <= 7'b1111101;
		7: SEG[6:0] <= 7'b0000111;
		8: SEG[6:0] <= 7'b1111111;
		9: SEG[6:0] <= 7'b1101111;
		10: SEG[6:0] <= 7'b1110111;
		11: SEG[6:0] <= 7'b1111100;
		12: SEG[6:0] <= 7'b0111001;
		13: SEG[6:0] <= 7'b1011110;
		14: SEG[6:0] <= 7'b1111001;
		15: SEG[6:0] <= 7'b1110001;

		// Letras e Símbolos

		16: SEG[6:0] <= 7'b1110111;
		17: SEG[6:0] <= 7'b1111100;
		18: SEG[6:0] <= 7'b0111001;
		19: SEG[6:0] <= 7'b1011000;
		20: SEG[6:0] <= 7'b1011110;
		21: SEG[6:0] <= 7'b1111001;
		22: SEG[6:0] <= 7'b1110001;
		23: SEG[6:0] <= 7'b1101111;
		24: SEG[6:0] <= 7'b1110110;
		25: SEG[6:0] <= 7'b1110100;
		26: SEG[6:0] <= 7'b0000100;
		27: SEG[6:0] <= 7'b0000110;
		28: SEG[6:0] <= 7'b0011110;
		29: SEG[6:0] <= 7'b0111000;
		30: SEG[6:0] <= 7'b1010100;
		31: SEG[6:0] <= 7'b0111111;
		32: SEG[6:0] <= 7'b1011100;
		33: SEG[6:0] <= 7'b1110011;
		34: SEG[6:0] <= 7'b1100111;
		35: SEG[6:0] <= 7'b1010000;
		36: SEG[6:0] <= 7'b1101101;
		37: SEG[6:0] <= 7'b1111000;
		38: SEG[6:0] <= 7'b0111110;
		39: SEG[6:0] <= 7'b0011100;
		40: SEG[6:0] <= 7'b1101110;
		41: SEG[6:0] <= 7'b1100011;

	default:
		SEG[6:0] <= 7'b1000000;
	endcase
end